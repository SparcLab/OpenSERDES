* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599667004215
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599667004212
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Inverter0 GND VDD INP OUT
** N=46 EP=4 IP=8 FDC=4
M0 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3140 $Y=1490 $D=9
M1 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2915 $Y=7755 $D=79
M2 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3345 $Y=7755 $D=79
X3 GND VDD Dpar a=11.524 p=15.02 m=1 $[nwdiode] $X=1790 $Y=7575 $D=191
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599667004219
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_CDNS_599667004217 2 3 4
** N=24 EP=3 IP=6 FDC=1
*.SEEDPROM
M0 4 3 2 2 pshort L=0.15 W=7 m=1 r=46.6667 a=1.05 p=14.3 mult=1 $X=0 $Y=0 $D=79
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_5996670042112
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_CDNS_5996670042110 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 4 2 3 1 nshort L=0.15 W=7 m=1 r=46.6667 a=1.05 p=14.3 mult=1 $X=0 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT NAND GND INP1 INP2 VDD OUT
** N=44 EP=5 IP=16 FDC=6
X0 GND VDD Dpar a=12.6592 p=18.16 m=1 $[nwdiode] $X=2130 $Y=9720 $D=191
X1 GND VDD Dpar a=12.6592 p=18.16 m=1 $[nwdiode] $X=5305 $Y=9705 $D=191
X2 VDD INP1 OUT pfet_CDNS_599667004217 $T=3255 9900 0 0 $X=2130 $Y=9720
X3 VDD INP2 OUT pfet_CDNS_599667004217 $T=6430 9885 0 0 $X=5305 $Y=9705
X4 GND INP1 6 OUT nfet_CDNS_5996670042110 $T=3255 1885 0 0 $X=2865 $Y=1755
X5 GND INP2 GND 6 nfet_CDNS_5996670042110 $T=6580 1885 1 180 $X=6040 $Y=1755
.ENDS
***************************************
.SUBCKT DFF GND D CLK Q_BAR Q VDD
** N=14 EP=6 IP=48 FDC=56
X0 GND VDD D 3 Inverter0 $T=1190 11745 0 0 $X=2375 $Y=12455
X1 GND VDD CLK 7 Inverter0 $T=27430 11745 0 0 $X=28615 $Y=12455
X2 GND D CLK VDD 12 NAND $T=5030 18685 0 0 $X=6420 $Y=19170
X3 GND 3 CLK VDD 11 NAND $T=5035 685 0 0 $X=6425 $Y=1170
X4 GND 11 6 VDD 5 NAND $T=12575 830 0 0 $X=13965 $Y=1315
X5 GND 12 5 VDD 6 NAND $T=12685 18715 0 0 $X=14075 $Y=19200
X6 GND 5 7 VDD 13 NAND $T=20810 830 0 0 $X=22200 $Y=1315
X7 GND 6 7 VDD 14 NAND $T=20920 18715 0 0 $X=22310 $Y=19200
X8 GND 13 Q VDD Q_BAR NAND $T=31545 830 0 0 $X=32935 $Y=1315
X9 GND 14 Q_BAR VDD Q NAND $T=31655 18715 0 0 $X=33045 $Y=19200
.ENDS
***************************************
