* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_3 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=0.59 W=0.55 m=1 r=0.932203 a=0.3245 p=2.28 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=0.59 W=0.87 m=1 r=1.47458 a=0.5133 p=2.92 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 5440 1 0 $X=-190 $Y=2480
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=4 FDC=8
*.SEEDPROM
X0 1 2 ICV_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_1 $T=0 5440 0 0 $X=-190 $Y=5200
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=4 FDC=16
*.SEEDPROM
X0 1 2 ICV_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_2 $T=0 10880 0 0 $X=-190 $Y=10640
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.05 W=0.55 m=1 r=0.52381 a=0.5775 p=3.2 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.05 W=0.87 m=1 r=0.828571 a=0.9135 p=3.84 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_6 VNB VPB VGND VPWR
** N=14 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.97 W=0.55 m=1 r=0.279188 a=1.0835 p=5.04 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.97 W=0.87 m=1 r=0.441624 a=1.7139 p=5.68 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_8 VNB VPB VGND VPWR
** N=16 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=2.89 W=0.55 m=1 r=0.190311 a=1.5895 p=6.88 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=2.89 W=0.87 m=1 r=0.301038 a=2.5143 p=7.52 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_5 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5060 0 1 180 $X=3490 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__buf_1 VNB VPB A VPWR X VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND A 7 VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 X 7 VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR A 7 VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 X 7 VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__diode_2 VNB DIODE
** N=9 EP=2 IP=0 FDC=1
*.SEEDPROM
D0 VNB DIODE ndiode AREA=0.4347 PJ=2.64 m=1 ahftempperim=2.64 $X=155 $Y=195 $D=167
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_7 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_8 1 2
** N=2 EP=2 IP=4 FDC=4
*.SEEDPROM
X1 1 2 ICV_7 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_12 VNB VPB VGND VPWR
** N=18 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=4.73 W=0.55 m=1 r=0.116279 a=2.6015 p=10.56 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=4.73 W=0.87 m=1 r=0.183932 a=4.1151 p=11.2 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_11 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_12 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor2_4 VNB VPB A B VPWR Y VGND
** N=51 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M9 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M10 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M11 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M12 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M13 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M14 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M15 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__inv_8 VNB VPB A VPWR Y VGND
** N=48 EP=6 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=560 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=980 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1400 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1820 $Y=235 $D=9
M4 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2240 $Y=235 $D=9
M5 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2660 $Y=235 $D=9
M6 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3080 $Y=235 $D=9
M7 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3500 $Y=235 $D=9
M8 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=560 $Y=1485 $D=89
M9 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=980 $Y=1485 $D=89
M10 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1400 $Y=1485 $D=89
M11 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1820 $Y=1485 $D=89
M12 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2240 $Y=1485 $D=89
M13 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2660 $Y=1485 $D=89
M14 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3080 $Y=1485 $D=89
M15 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3500 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4
** N=4 EP=4 IP=10 FDC=18
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 4 2 3 1 sky130_fd_sc_hd__inv_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_14 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3
** N=3 EP=3 IP=5 FDC=3
*.SEEDPROM
X1 1 2 3 ICV_15 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_17 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_18 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_7 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 ICV_18 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_21 1 3 4
** N=4 EP=3 IP=10 FDC=2
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 4 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_24 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21oi_4 VNB VPB B1 A2 A1 Y VPWR VGND
** N=57 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2590 $Y=235 $D=9
M6 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3020 $Y=235 $D=9
M7 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3450 $Y=235 $D=9
M8 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3880 $Y=235 $D=9
M9 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4310 $Y=235 $D=9
M10 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4740 $Y=235 $D=9
M11 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5170 $Y=235 $D=9
M12 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M13 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M14 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M15 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M16 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2150 $Y=1485 $D=89
M17 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2590 $Y=1485 $D=89
M18 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3020 $Y=1485 $D=89
M19 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3450 $Y=1485 $D=89
M20 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3880 $Y=1485 $D=89
M21 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4310 $Y=1485 $D=89
M22 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4740 $Y=1485 $D=89
M23 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor3_4 VNB VPB A B C VPWR Y VGND
** N=63 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3775 $Y=235 $D=9
M9 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4195 $Y=235 $D=9
M10 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4615 $Y=235 $D=9
M11 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5035 $Y=235 $D=9
M12 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M13 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M14 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M15 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M16 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M17 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M18 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M19 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
M20 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3775 $Y=1485 $D=89
M21 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4195 $Y=1485 $D=89
M22 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4615 $Y=1485 $D=89
M23 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5035 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4
** N=4 EP=4 IP=10 FDC=18
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 4 2 3 1 sky130_fd_sc_hd__inv_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3
** N=3 EP=3 IP=7 FDC=5
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 3 ICV_9 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o22a_4 VNB VPB B1 B2 A1 A2 VPWR X VGND
** N=65 EP=9 IP=0 FDC=24
*.SEEDPROM
M0 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=480 $Y=235 $D=9
M1 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=900 $Y=235 $D=9
M2 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=9
M3 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1740 $Y=235 $D=9
M4 10 B1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2680 $Y=235 $D=9
M5 13 B2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3100 $Y=235 $D=9
M6 10 B2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3520 $Y=235 $D=9
M7 13 B1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3940 $Y=235 $D=9
M8 VGND A1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4440 $Y=235 $D=9
M9 13 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4860 $Y=235 $D=9
M10 VGND A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5280 $Y=235 $D=9
M11 13 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5700 $Y=235 $D=9
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=480 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=900 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M16 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2680 $Y=1485 $D=89
M17 10 B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3100 $Y=1485 $D=89
M18 11 B2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3520 $Y=1485 $D=89
M19 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3940 $Y=1485 $D=89
M20 12 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4440 $Y=1485 $D=89
M21 10 A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4860 $Y=1485 $D=89
M22 12 A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5280 $Y=1485 $D=89
M23 VPWR A1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5700 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=17
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 2 4 1 sky130_fd_sc_hd__inv_8 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nand2_4 VNB VPB B A VPWR Y VGND
** N=50 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 8 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 Y A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 8 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M9 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M10 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M11 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M12 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M13 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M14 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M15 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a2bb2o_4 VNB VPB B1 B2 A1_N A2_N VPWR X VGND
** N=75 EP=9 IP=0 FDC=28
*.SEEDPROM
M0 14 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 11 B2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 14 B2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 VGND B1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 11 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 VGND 10 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 10 A1_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3435 $Y=235 $D=9
M7 VGND A2_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3855 $Y=235 $D=9
M8 10 A2_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 VGND A1_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5115 $Y=235 $D=9
M11 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5535 $Y=235 $D=9
M12 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5955 $Y=235 $D=9
M13 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6375 $Y=235 $D=9
M14 VPWR B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M15 12 B2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M16 VPWR B2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M17 12 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M18 11 10 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M19 12 10 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M20 13 A1_N VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3435 $Y=1485 $D=89
M21 10 A2_N 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3855 $Y=1485 $D=89
M22 13 A2_N 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4275 $Y=1485 $D=89
M23 VPWR A1_N 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4695 $Y=1485 $D=89
M24 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5115 $Y=1485 $D=89
M25 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5535 $Y=1485 $D=89
M26 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5955 $Y=1485 $D=89
M27 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6375 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_21 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_21 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3
** N=3 EP=3 IP=7 FDC=5
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 3 ICV_9 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and2_4 VNB VPB A B VPWR X VGND
** N=38 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 9 A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=760 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1335 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1765 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2195 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2625 $Y=235 $D=9
M6 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M7 VPWR B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1335 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1765 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2195 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2625 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or2_4 VNB VPB B A VPWR X VGND
** N=37 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1740 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2580 $Y=235 $D=9
M6 9 B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=455 $Y=1485 $D=89
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2160 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4_4 VNB VPB A B C D VPWR X VGND
** N=44 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 11 A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 12 B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=790 $Y=235 $D=8
M2 13 C 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1275 $Y=235 $D=8
M3 VGND D 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1860 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2335 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2755 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3175 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3595 $Y=235 $D=9
M8 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M9 VPWR B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M10 10 C VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1275 $Y=1485 $D=89
M11 VPWR D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1855 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2335 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2755 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3175 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3595 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_15 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 4 5 ICV_21 $T=3220 0 0 0 $X=3030 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
** N=109 EP=9 IP=0 FDC=40
*.SEEDPROM
M0 13 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND B1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 13 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 Y B2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 13 B2 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 Y B2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 13 B2 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 VGND B1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 Y 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3755 $Y=235 $D=9
M9 VGND 10 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4175 $Y=235 $D=9
M10 Y 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4595 $Y=235 $D=9
M11 VGND 10 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5015 $Y=235 $D=9
M12 10 A1_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5955 $Y=235 $D=9
M13 VGND A1_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6375 $Y=235 $D=9
M14 10 A1_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6795 $Y=235 $D=9
M15 VGND A1_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7215 $Y=235 $D=9
M16 10 A2_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7635 $Y=235 $D=9
M17 VGND A2_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8055 $Y=235 $D=9
M18 10 A2_N VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8475 $Y=235 $D=9
M19 VGND A2_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8895 $Y=235 $D=9
M20 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M21 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M22 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M23 11 B2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M24 VPWR B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M25 11 B2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M26 VPWR B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M27 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
M28 Y 10 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3755 $Y=1485 $D=89
M29 11 10 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4175 $Y=1485 $D=89
M30 Y 10 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4595 $Y=1485 $D=89
M31 11 10 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5015 $Y=1485 $D=89
M32 VPWR A1_N 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5955 $Y=1485 $D=89
M33 12 A1_N VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6375 $Y=1485 $D=89
M34 VPWR A1_N 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6795 $Y=1485 $D=89
M35 12 A1_N VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7215 $Y=1485 $D=89
M36 10 A2_N 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7635 $Y=1485 $D=89
M37 12 A2_N 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8055 $Y=1485 $D=89
M38 10 A2_N 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8475 $Y=1485 $D=89
M39 12 A2_N 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8895 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dfrtp_4 VNB VPB CLK D RESET_B VPWR Q VGND
** N=88 EP=8 IP=0 FDC=34
*.SEEDPROM
M0 VGND CLK 9 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 10 9 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 15 D VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2090 $Y=235 $D=9
M3 12 9 15 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=2565 $Y=235 $D=9
M4 18 10 12 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=3045 $Y=235 $D=9
M5 19 11 18 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3875 $Y=235 $D=8
M6 VGND RESET_B 19 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4235 $Y=235 $D=9
M7 11 12 VGND VNB nshort L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=4895 $Y=235 $D=9
M8 14 10 11 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5390 $Y=235 $D=9
M9 20 9 14 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5935 $Y=235 $D=9
M10 VGND 13 20 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M11 21 RESET_B VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=235 $D=9
M12 13 14 21 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7615 $Y=235 $D=9
M13 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8555 $Y=235 $D=9
M14 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8975 $Y=235 $D=9
M15 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9395 $Y=235 $D=9
M16 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9815 $Y=235 $D=9
M17 VPWR CLK 9 VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M18 10 9 VPWR VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M19 15 D VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2150 $Y=2065 $D=89
M20 12 10 15 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2610 $Y=2065 $D=89
M21 16 9 12 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3105 $Y=2065 $D=89
M22 VPWR 11 16 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3805 $Y=2065 $D=89
M23 16 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4290 $Y=2065 $D=89
M24 11 12 VPWR VPB phighvt L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=5275 $Y=1645 $D=89
M25 14 9 11 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5770 $Y=2065 $D=89
M26 17 10 14 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6200 $Y=2065 $D=89
M27 VPWR 13 17 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6620 $Y=2065 $D=89
M28 13 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=2065 $D=89
M29 VPWR 14 13 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7580 $Y=2065 $D=89
M30 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8555 $Y=1485 $D=89
M31 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8975 $Y=1485 $D=89
M32 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9395 $Y=1485 $D=89
M33 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9815 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=13
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__and2_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_35 1 3 4 5
** N=5 EP=4 IP=9 FDC=3
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 4 5 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a211o_4 VNB VPB B1 C1 A2 A1 VPWR X VGND
** N=59 EP=9 IP=0 FDC=24
*.SEEDPROM
M0 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=790 $Y=235 $D=9
M1 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1220 $Y=235 $D=9
M2 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1650 $Y=235 $D=9
M3 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M4 10 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2530 $Y=235 $D=9
M5 VGND C1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3000 $Y=235 $D=9
M6 10 C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3485 $Y=235 $D=9
M7 VGND B1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4025 $Y=235 $D=9
M8 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4605 $Y=235 $D=9
M9 10 A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5035 $Y=235 $D=9
M10 15 A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5465 $Y=235 $D=9
M11 VGND A2 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5895 $Y=235 $D=9
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=825 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1685 $Y=1485 $D=89
M16 12 B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2625 $Y=1485 $D=89
M17 10 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3055 $Y=1485 $D=89
M18 13 C1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3485 $Y=1485 $D=89
M19 11 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3955 $Y=1485 $D=89
M20 VPWR A2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4495 $Y=1485 $D=89
M21 11 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5035 $Y=1485 $D=89
M22 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5465 $Y=1485 $D=89
M23 11 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5895 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4
** N=4 EP=4 IP=10 FDC=6
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=1380 0 0 0 $X=1190 $Y=-240
X1 1 2 3 2 4 1 sky130_fd_sc_hd__buf_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_39 1 3 4 5 6
** N=6 EP=5 IP=8 FDC=4
*.SEEDPROM
X0 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 5 6 ICV_21 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_9 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 4 5 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=15
*.SEEDPROM
X0 1 2 3 ICV_6 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__or2_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_42 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_43 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_15 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 4 5 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_44 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_21 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o21ai_4 VNB VPB A1 A2 B1 VPWR Y VGND
** N=52 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 VGND A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=425 $Y=235 $D=9
M1 10 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=855 $Y=235 $D=9
M2 VGND A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1285 $Y=235 $D=9
M3 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1715 $Y=235 $D=9
M4 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2145 $Y=235 $D=9
M5 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2575 $Y=235 $D=9
M6 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3005 $Y=235 $D=9
M7 10 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3475 $Y=235 $D=9
M8 Y B1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3905 $Y=235 $D=9
M9 10 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4335 $Y=235 $D=9
M10 Y B1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4765 $Y=235 $D=9
M11 10 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5195 $Y=235 $D=9
M12 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=425 $Y=1485 $D=89
M13 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=855 $Y=1485 $D=89
M14 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1285 $Y=1485 $D=89
M15 Y A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1715 $Y=1485 $D=89
M16 9 A2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2145 $Y=1485 $D=89
M17 Y A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2575 $Y=1485 $D=89
M18 9 A2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3005 $Y=1485 $D=89
M19 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3435 $Y=1485 $D=89
M20 Y B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3905 $Y=1485 $D=89
M21 VPWR B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4335 $Y=1485 $D=89
M22 Y B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4765 $Y=1485 $D=89
M23 VPWR B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5195 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_45 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_46 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_21 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=19
*.SEEDPROM
X0 1 2 4 2 3 1 sky130_fd_sc_hd__inv_8 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 2 5 ICV_33 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o21a_4 VNB VPB B1 A1 A2 VPWR X VGND
** N=53 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 9 B1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2640 $Y=235 $D=9
M5 12 B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3070 $Y=235 $D=9
M6 VGND A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M7 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4090 $Y=235 $D=9
M8 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4520 $Y=235 $D=9
M9 12 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4950 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=720 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1150 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1580 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2010 $Y=1485 $D=89
M14 9 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2460 $Y=1485 $D=89
M15 VPWR B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2890 $Y=1485 $D=89
M16 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3660 $Y=1485 $D=89
M17 9 A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4090 $Y=1485 $D=89
M18 11 A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4520 $Y=1485 $D=89
M19 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4950 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_50 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_51 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_52 1 3
** N=3 EP=2 IP=7 FDC=1
*.SEEDPROM
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_53 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_54 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_55 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_56 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X1 1 2 3 2 4 1 sky130_fd_sc_hd__buf_1 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_57 1 2 3 4
** N=4 EP=4 IP=8 FDC=16
*.SEEDPROM
X1 1 2 4 2 3 1 sky130_fd_sc_hd__inv_8 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_58 1 3 4
** N=4 EP=3 IP=6 FDC=2
*.SEEDPROM
X1 1 3 4 ICV_21 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_59 1 2 3 4
** N=4 EP=4 IP=6 FDC=4
*.SEEDPROM
X0 1 3 4 ICV_21 $T=1840 0 0 0 $X=1650 $Y=-240
X1 1 2 ICV_54 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_60 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__or2_4 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_61 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=3220 0 0 0 $X=3030 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__or2_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or4_4 VNB VPB D C B A VPWR X VGND
** N=46 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 10 D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND C 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=950 $Y=235 $D=9
M2 10 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1370 $Y=235 $D=9
M3 VGND A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1790 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2320 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2740 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3160 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M8 11 D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M9 12 C 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=950 $Y=1485 $D=88
M10 13 B 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1370 $Y=1485 $D=88
M11 VPWR A 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1790 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2320 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2740 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3160 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_62 1 3
** N=3 EP=2 IP=7 FDC=1
*.SEEDPROM
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_63 1 2 3
** N=3 EP=3 IP=7 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=2300 0 0 0 $X=2110 $Y=-240
X1 1 3 ICV_62 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21o_4 VNB VPB B1 A2 A1 VPWR X VGND
** N=55 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=850 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1280 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1710 $Y=235 $D=9
M4 9 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2675 $Y=235 $D=9
M5 VGND B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3095 $Y=235 $D=9
M6 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3555 $Y=235 $D=9
M7 9 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3935 $Y=235 $D=9
M8 12 A1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4355 $Y=235 $D=9
M9 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4775 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=850 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1280 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1710 $Y=1485 $D=89
M14 9 B1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2675 $Y=1485 $D=89
M15 10 B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3095 $Y=1485 $D=89
M16 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3515 $Y=1485 $D=89
M17 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3935 $Y=1485 $D=89
M18 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4355 $Y=1485 $D=89
M19 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4775 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 ICV_36 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_65 1 3 4
** N=4 EP=3 IP=6 FDC=2
*.SEEDPROM
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_66 1 2 3
** N=3 EP=3 IP=5 FDC=3
*.SEEDPROM
X1 1 2 3 ICV_33 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_67 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_15 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 4 5 ICV_21 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a32o_4 VNB VPB A3 A2 A1 B1 B2 VPWR X VGND
** N=67 EP=10 IP=0 FDC=28
*.SEEDPROM
M0 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 13 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 VGND A3 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 13 A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3435 $Y=235 $D=9
M7 14 A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3855 $Y=235 $D=9
M8 11 A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 14 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 11 B1 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5970 $Y=235 $D=9
M11 15 B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6390 $Y=235 $D=9
M12 VGND B2 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6855 $Y=235 $D=9
M13 15 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7275 $Y=235 $D=9
M14 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M15 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M16 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M17 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M18 12 A3 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M19 VPWR A3 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M20 VPWR A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3435 $Y=1485 $D=89
M21 12 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3855 $Y=1485 $D=89
M22 VPWR A1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4275 $Y=1485 $D=89
M23 12 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4695 $Y=1485 $D=89
M24 11 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6015 $Y=1485 $D=89
M25 12 B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6435 $Y=1485 $D=89
M26 11 B2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6855 $Y=1485 $D=89
M27 12 B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_68 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 ICV_33 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_70 1 2 3
** N=3 EP=3 IP=7 FDC=5
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=2300 0 0 0 $X=2110 $Y=-240
X1 1 2 3 ICV_36 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_71 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=13
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__or2_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_72 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=15
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__or2_4 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 2 6 ICV_33 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_73 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=5
*.SEEDPROM
X0 1 2 3 2 4 1 sky130_fd_sc_hd__buf_1 $T=1840 0 0 0 $X=1650 $Y=-240
X1 1 5 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a2111oi_4 VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
** N=104 EP=10 IP=0 FDC=40
*.SEEDPROM
M0 Y D1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND D1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y D1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1265 $Y=235 $D=9
M3 VGND D1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1695 $Y=235 $D=9
M4 Y C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2205 $Y=235 $D=9
M5 VGND C1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2635 $Y=235 $D=9
M6 Y C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3065 $Y=235 $D=9
M7 VGND C1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3495 $Y=235 $D=9
M8 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4035 $Y=235 $D=9
M9 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4465 $Y=235 $D=9
M10 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4895 $Y=235 $D=9
M11 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5325 $Y=235 $D=9
M12 Y A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6305 $Y=235 $D=9
M13 14 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6735 $Y=235 $D=9
M14 Y A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7165 $Y=235 $D=9
M15 14 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7595 $Y=235 $D=9
M16 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8120 $Y=235 $D=9
M17 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8550 $Y=235 $D=9
M18 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8980 $Y=235 $D=9
M19 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9410 $Y=235 $D=9
M20 Y D1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=405 $Y=1485 $D=89
M21 11 D1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M22 Y D1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1265 $Y=1485 $D=89
M23 11 D1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1695 $Y=1485 $D=89
M24 12 C1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2125 $Y=1485 $D=89
M25 11 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2555 $Y=1485 $D=89
M26 12 C1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2985 $Y=1485 $D=89
M27 11 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3415 $Y=1485 $D=89
M28 12 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4365 $Y=1485 $D=89
M29 13 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4795 $Y=1485 $D=89
M30 12 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5225 $Y=1485 $D=89
M31 13 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5655 $Y=1485 $D=89
M32 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6095 $Y=1485 $D=89
M33 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6525 $Y=1485 $D=89
M34 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6955 $Y=1485 $D=89
M35 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7405 $Y=1485 $D=89
M36 VPWR A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7955 $Y=1485 $D=89
M37 13 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8385 $Y=1485 $D=89
M38 VPWR A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8905 $Y=1485 $D=89
M39 13 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9335 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_74 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a22oi_4 VNB VPB B2 B1 A1 A2 Y VPWR VGND
** N=94 EP=9 IP=0 FDC=32
*.SEEDPROM
M0 VGND B2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 11 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND B2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 11 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 11 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 Y B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 11 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 Y A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 12 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 Y A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5115 $Y=235 $D=9
M11 12 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5535 $Y=235 $D=9
M12 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5955 $Y=235 $D=9
M13 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6375 $Y=235 $D=9
M14 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6795 $Y=235 $D=9
M15 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7215 $Y=235 $D=9
M16 Y B2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M17 10 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M18 Y B2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M19 10 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M20 Y B1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M21 10 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M22 Y B1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M23 10 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
M24 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4275 $Y=1485 $D=89
M25 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4695 $Y=1485 $D=89
M26 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5115 $Y=1485 $D=89
M27 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5535 $Y=1485 $D=89
M28 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5955 $Y=1485 $D=89
M29 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6375 $Y=1485 $D=89
M30 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6795 $Y=1485 $D=89
M31 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7215 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_75 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_76 1 3 4 5
** N=5 EP=4 IP=7 FDC=3
*.SEEDPROM
X0 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 5 ICV_62 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dfstp_4 VNB VPB CLK D SET_B VPWR Q VGND
** N=94 EP=8 IP=0 FDC=40
*.SEEDPROM
M0 VGND CLK 9 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 10 9 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 16 D VGND VNB nshort L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=1755 $Y=235 $D=9
M3 12 9 16 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=2230 $Y=235 $D=9
M4 20 10 12 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=2780 $Y=235 $D=9
M5 VGND 11 20 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3260 $Y=235 $D=9
M6 21 SET_B VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3830 $Y=235 $D=9
M7 11 12 21 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4190 $Y=235 $D=9
M8 22 12 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5130 $Y=235 $D=9
M9 14 10 22 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5490 $Y=235 $D=9
M10 23 9 14 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5970 $Y=235 $D=9
M11 24 13 23 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6330 $Y=235 $D=8
M12 VGND SET_B 24 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6690 $Y=235 $D=9
M13 13 14 VGND VNB nshort L=0.15 W=0.54 m=1 r=3.6 a=0.081 p=1.38 mult=1 $X=7310 $Y=235 $D=9
M14 VGND 14 15 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8250 $Y=235 $D=9
M15 Q 15 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8725 $Y=235 $D=9
M16 VGND 15 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9145 $Y=235 $D=9
M17 Q 15 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9565 $Y=235 $D=9
M18 VGND 15 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9985 $Y=235 $D=9
M19 Q 15 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=10405 $Y=235 $D=9
M20 VPWR CLK 9 VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M21 10 9 VPWR VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M22 16 D VPWR VPB phighvt L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=1755 $Y=1645 $D=89
M23 12 10 16 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2240 $Y=2065 $D=89
M24 17 9 12 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2660 $Y=2065 $D=89
M25 VPWR 11 17 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3260 $Y=2065 $D=89
M26 11 SET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3790 $Y=2065 $D=89
M27 VPWR 12 11 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4210 $Y=2065 $D=89
M28 18 12 VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4630 $Y=2065 $D=89
M29 14 9 18 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4990 $Y=2065 $D=89
M30 19 10 14 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5530 $Y=2065 $D=89
M31 VPWR 13 19 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5890 $Y=2065 $D=89
M32 VPWR SET_B 14 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6830 $Y=2065 $D=89
M33 13 14 VPWR VPB phighvt L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=7310 $Y=1645 $D=89
M34 VPWR 14 15 VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=8250 $Y=1845 $D=89
M35 Q 15 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8725 $Y=1485 $D=89
M36 VPWR 15 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9145 $Y=1485 $D=89
M37 Q 15 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9565 $Y=1485 $D=89
M38 VPWR 15 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9985 $Y=1485 $D=89
M39 Q 15 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=10405 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a32oi_4 VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
** N=96 EP=10 IP=0 FDC=40
*.SEEDPROM
M0 VGND B2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 12 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND B2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 12 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y B1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 12 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 Y B1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 12 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 Y A1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 13 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 Y A1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5115 $Y=235 $D=9
M11 13 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5535 $Y=235 $D=9
M12 14 A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6095 $Y=235 $D=9
M13 13 A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6515 $Y=235 $D=9
M14 14 A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6935 $Y=235 $D=9
M15 13 A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7355 $Y=235 $D=9
M16 14 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8295 $Y=235 $D=9
M17 VGND A3 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8715 $Y=235 $D=9
M18 14 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9135 $Y=235 $D=9
M19 VGND A3 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9555 $Y=235 $D=9
M20 Y B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M21 11 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M22 Y B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M23 11 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M24 Y B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M25 11 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M26 Y B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M27 11 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
M28 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3775 $Y=1485 $D=89
M29 11 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4195 $Y=1485 $D=89
M30 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4615 $Y=1485 $D=89
M31 11 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5440 $Y=1485 $D=89
M32 VPWR A2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6095 $Y=1485 $D=89
M33 11 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6515 $Y=1485 $D=89
M34 VPWR A2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6935 $Y=1485 $D=89
M35 11 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7355 $Y=1485 $D=89
M36 VPWR A3 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8295 $Y=1485 $D=89
M37 11 A3 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8715 $Y=1485 $D=89
M38 VPWR A3 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9135 $Y=1485 $D=89
M39 11 A3 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9555 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or3_4 VNB VPB C B A VPWR X VGND
** N=49 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 VGND C 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 9 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2185 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2605 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3025 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3445 $Y=235 $D=9
M7 10 C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M8 11 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=88
M9 VPWR A 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2185 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2605 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3025 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3445 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_77 1 2 3
** N=3 EP=3 IP=7 FDC=5
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 3 ICV_9 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_78 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=14
*.SEEDPROM
X0 1 3 4 ICV_21 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 5 6 2 7 1 sky130_fd_sc_hd__and2_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_79 1 2 3
** N=3 EP=3 IP=7 FDC=5
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 3 ICV_9 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_80 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o41a_4 VNB VPB B1 A4 A3 A2 A1 VPWR X VGND
** N=92 EP=10 IP=0 FDC=28
*.SEEDPROM
M0 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 11 B1 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2595 $Y=235 $D=9
M5 15 B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3015 $Y=235 $D=9
M6 VGND A4 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3455 $Y=235 $D=9
M7 15 A4 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3875 $Y=235 $D=9
M8 VGND A3 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4295 $Y=235 $D=9
M9 15 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4715 $Y=235 $D=9
M10 VGND A2 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5155 $Y=235 $D=9
M11 15 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5915 $Y=235 $D=9
M12 VGND A1 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6535 $Y=235 $D=9
M13 15 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6955 $Y=235 $D=9
M14 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M15 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M16 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M17 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M18 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M19 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M20 11 A4 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3455 $Y=1485 $D=89
M21 12 A4 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3875 $Y=1485 $D=89
M22 13 A3 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4295 $Y=1485 $D=89
M23 12 A3 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4715 $Y=1485 $D=89
M24 13 A2 14 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5695 $Y=1485 $D=89
M25 14 A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6115 $Y=1485 $D=89
M26 VPWR A1 14 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6535 $Y=1485 $D=89
M27 14 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6955 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor4_4 VNB VPB A B C D VPWR Y VGND
** N=94 EP=9 IP=0 FDC=32
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4295 $Y=235 $D=9
M9 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4715 $Y=235 $D=9
M10 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5135 $Y=235 $D=9
M11 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5555 $Y=235 $D=9
M12 Y D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5975 $Y=235 $D=9
M13 VGND D Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6395 $Y=235 $D=9
M14 Y D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6815 $Y=235 $D=9
M15 VGND D Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7235 $Y=235 $D=9
M16 VPWR A 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M17 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M18 VPWR A 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M19 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M20 11 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M21 10 B 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M22 11 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M23 10 B 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
M24 11 C 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4295 $Y=1485 $D=89
M25 12 C 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4715 $Y=1485 $D=89
M26 11 C 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5135 $Y=1485 $D=89
M27 12 C 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5555 $Y=1485 $D=89
M28 Y D 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5975 $Y=1485 $D=89
M29 12 D Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6395 $Y=1485 $D=89
M30 Y D 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6815 $Y=1485 $D=89
M31 12 D Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7235 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_81 1 2 3
** N=3 EP=3 IP=5 FDC=5
*.SEEDPROM
X0 1 2 ICV_4 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 2 3 ICV_15 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_82 1 2 3
** N=3 EP=3 IP=5 FDC=3
*.SEEDPROM
X1 1 2 3 ICV_36 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and3_4 VNB VPB A B C VPWR X VGND
** N=43 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 10 A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=775 $Y=235 $D=9
M1 11 B 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=8
M2 VGND C 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1680 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2255 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2685 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3115 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3545 $Y=235 $D=9
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=775 $Y=1485 $D=89
M8 9 B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1750 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2255 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2685 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3115 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3545 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_83 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 3 4 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 ICV_37 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o32ai_4 VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
** N=112 EP=10 IP=0 FDC=40
*.SEEDPROM
M0 Y B2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 14 B2 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 Y B2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 14 B2 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y B1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2090 $Y=235 $D=9
M5 14 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2510 $Y=235 $D=9
M6 Y B1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2930 $Y=235 $D=9
M7 14 B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3350 $Y=235 $D=9
M8 VGND A3 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3770 $Y=235 $D=9
M9 14 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4190 $Y=235 $D=9
M10 VGND A3 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4610 $Y=235 $D=9
M11 14 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5190 $Y=235 $D=9
M12 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5970 $Y=235 $D=9
M13 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6390 $Y=235 $D=9
M14 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6810 $Y=235 $D=9
M15 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7230 $Y=235 $D=9
M16 VGND A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8170 $Y=235 $D=9
M17 14 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8590 $Y=235 $D=9
M18 VGND A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9010 $Y=235 $D=9
M19 14 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9525 $Y=235 $D=9
M20 Y B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M21 11 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M22 Y B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M23 11 B2 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M24 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2090 $Y=1485 $D=89
M25 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2510 $Y=1485 $D=89
M26 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2930 $Y=1485 $D=89
M27 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3350 $Y=1485 $D=89
M28 Y A3 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4290 $Y=1485 $D=89
M29 12 A3 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4710 $Y=1485 $D=89
M30 Y A3 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5130 $Y=1485 $D=89
M31 12 A3 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5550 $Y=1485 $D=89
M32 13 A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5970 $Y=1485 $D=89
M33 12 A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6390 $Y=1485 $D=89
M34 13 A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6810 $Y=1485 $D=89
M35 12 A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7230 $Y=1485 $D=89
M36 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8170 $Y=1485 $D=89
M37 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8590 $Y=1485 $D=89
M38 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9010 $Y=1485 $D=89
M39 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9525 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_84 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_6 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 4 5 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_85 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=15
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_4 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 2 6 ICV_33 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_86 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=15
*.SEEDPROM
X0 1 2 3 ICV_15 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__or2_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21boi_4 VNB VPB B1_N A2 A1 VPWR Y VGND
** N=63 EP=8 IP=0 FDC=26
*.SEEDPROM
M0 VGND B1_N 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=550 $Y=235 $D=9
M1 Y 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1080 $Y=235 $D=9
M2 VGND 9 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1510 $Y=235 $D=9
M3 Y 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1940 $Y=235 $D=9
M4 VGND 9 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2370 $Y=235 $D=9
M5 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3140 $Y=235 $D=9
M6 Y A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3570 $Y=235 $D=9
M7 11 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4000 $Y=235 $D=9
M8 Y A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4430 $Y=235 $D=9
M9 11 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4860 $Y=235 $D=9
M10 VGND A2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5290 $Y=235 $D=9
M11 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5720 $Y=235 $D=9
M12 VGND A2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6150 $Y=235 $D=9
M13 VPWR B1_N 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=430 $Y=1485 $D=89
M14 Y 9 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1380 $Y=1485 $D=89
M15 10 9 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1810 $Y=1485 $D=89
M16 Y 9 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2240 $Y=1485 $D=89
M17 10 9 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2670 $Y=1485 $D=89
M18 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3130 $Y=1485 $D=89
M19 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3570 $Y=1485 $D=89
M20 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4000 $Y=1485 $D=89
M21 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4430 $Y=1485 $D=89
M22 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4860 $Y=1485 $D=89
M23 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5290 $Y=1485 $D=89
M24 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5720 $Y=1485 $D=89
M25 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6150 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_16 VNB VPB A VPWR X VGND
** N=79 EP=6 IP=0 FDC=40
*.SEEDPROM
M0 7 A VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=830 $Y=235 $D=9
M2 7 A VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1260 $Y=235 $D=9
M3 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1690 $Y=235 $D=9
M4 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2120 $Y=235 $D=9
M5 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2550 $Y=235 $D=9
M6 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2980 $Y=235 $D=9
M7 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3410 $Y=235 $D=9
M8 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3840 $Y=235 $D=9
M9 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4270 $Y=235 $D=9
M10 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4700 $Y=235 $D=9
M11 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5130 $Y=235 $D=9
M12 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5555 $Y=235 $D=9
M13 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5985 $Y=235 $D=9
M14 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M15 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6845 $Y=235 $D=9
M16 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7275 $Y=235 $D=9
M17 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7705 $Y=235 $D=9
M18 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8135 $Y=235 $D=9
M19 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8565 $Y=235 $D=9
M20 7 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M21 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M22 7 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M23 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M24 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2120 $Y=1485 $D=89
M25 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2550 $Y=1485 $D=89
M26 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2980 $Y=1485 $D=89
M27 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3410 $Y=1485 $D=89
M28 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3840 $Y=1485 $D=89
M29 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4270 $Y=1485 $D=89
M30 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4700 $Y=1485 $D=89
M31 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5130 $Y=1485 $D=89
M32 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5555 $Y=1485 $D=89
M33 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5985 $Y=1485 $D=89
M34 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6415 $Y=1485 $D=89
M35 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6845 $Y=1485 $D=89
M36 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
M37 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7705 $Y=1485 $D=89
M38 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8135 $Y=1485 $D=89
M39 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8565 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_87 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 2 3 ICV_20 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 4 5 ICV_21 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_88 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_14 $T=11040 0 0 0 $X=10850 $Y=-240
X1 1 2 ICV_42 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_89 1 2
** N=2 EP=2 IP=4 FDC=12
*.SEEDPROM
X0 1 2 ICV_88 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_88 $T=14260 0 0 0 $X=14070 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21bo_4 VNB VPB B1_N A2 A1 VPWR X VGND
** N=52 EP=8 IP=0 FDC=22
*.SEEDPROM
M0 VGND B1_N 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=595 $Y=235 $D=9
M1 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1025 $Y=235 $D=9
M2 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1455 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1885 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2315 $Y=235 $D=9
M5 9 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3275 $Y=235 $D=9
M6 VGND 10 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3695 $Y=235 $D=9
M7 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4155 $Y=235 $D=9
M8 9 A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4535 $Y=235 $D=9
M9 13 A1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4955 $Y=235 $D=9
M10 VGND A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5375 $Y=235 $D=9
M11 VPWR B1_N 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=595 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1025 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1455 $Y=1485 $D=89
M14 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1885 $Y=1485 $D=89
M15 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2315 $Y=1485 $D=89
M16 9 10 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3275 $Y=1485 $D=89
M17 11 10 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3695 $Y=1485 $D=89
M18 VPWR A2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4115 $Y=1485 $D=89
M19 11 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4535 $Y=1485 $D=89
M20 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4955 $Y=1485 $D=89
M21 11 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5375 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__xor2_4 VNB VPB A B VPWR X VGND
** N=100 EP=7 IP=0 FDC=40
*.SEEDPROM
M0 8 A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=410 $Y=235 $D=9
M1 VGND A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 8 A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1250 $Y=235 $D=9
M3 VGND A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1670 $Y=235 $D=9
M4 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2090 $Y=235 $D=9
M5 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2510 $Y=235 $D=9
M6 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2930 $Y=235 $D=9
M7 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3350 $Y=235 $D=9
M8 X B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4290 $Y=235 $D=9
M9 11 B X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4710 $Y=235 $D=9
M10 X B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5130 $Y=235 $D=9
M11 11 B X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5550 $Y=235 $D=9
M12 VGND A 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5970 $Y=235 $D=9
M13 11 A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6390 $Y=235 $D=9
M14 VGND A 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6810 $Y=235 $D=9
M15 11 A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7230 $Y=235 $D=9
M16 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8180 $Y=235 $D=9
M17 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8600 $Y=235 $D=9
M18 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9020 $Y=235 $D=9
M19 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9440 $Y=235 $D=9
M20 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=410 $Y=1485 $D=89
M21 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M22 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1250 $Y=1485 $D=89
M23 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1670 $Y=1485 $D=89
M24 8 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2090 $Y=1485 $D=89
M25 9 B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2510 $Y=1485 $D=89
M26 8 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2930 $Y=1485 $D=89
M27 9 B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3350 $Y=1485 $D=89
M28 VPWR B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4290 $Y=1485 $D=89
M29 10 B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4710 $Y=1485 $D=89
M30 VPWR B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5130 $Y=1485 $D=89
M31 10 B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5550 $Y=1485 $D=89
M32 VPWR A 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5970 $Y=1485 $D=89
M33 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6390 $Y=1485 $D=89
M34 VPWR A 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6810 $Y=1485 $D=89
M35 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7230 $Y=1485 $D=89
M36 10 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8180 $Y=1485 $D=89
M37 X 8 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8600 $Y=1485 $D=89
M38 10 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9020 $Y=1485 $D=89
M39 X 8 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9440 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a2111o_4 VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
** N=79 EP=10 IP=0 FDC=28
*.SEEDPROM
M0 VGND D1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=485 $Y=235 $D=9
M1 11 D1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=915 $Y=235 $D=9
M2 VGND C1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1345 $Y=235 $D=9
M3 11 C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1810 $Y=235 $D=9
M4 VGND B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2295 $Y=235 $D=9
M5 11 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3265 $Y=235 $D=9
M6 15 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3700 $Y=235 $D=9
M7 11 A1 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4130 $Y=235 $D=9
M8 15 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5110 $Y=235 $D=9
M9 VGND A2 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5540 $Y=235 $D=9
M10 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5970 $Y=235 $D=9
M11 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6400 $Y=235 $D=9
M12 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6830 $Y=235 $D=9
M13 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7260 $Y=235 $D=9
M14 11 D1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M15 12 D1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=845 $Y=1485 $D=89
M16 13 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1275 $Y=1485 $D=89
M17 12 C1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1705 $Y=1485 $D=89
M18 13 B1 14 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2645 $Y=1485 $D=89
M19 14 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3075 $Y=1485 $D=89
M20 VPWR A1 14 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3740 $Y=1485 $D=89
M21 14 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4170 $Y=1485 $D=89
M22 14 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5110 $Y=1485 $D=89
M23 VPWR A2 14 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5540 $Y=1485 $D=89
M24 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5970 $Y=1485 $D=89
M25 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6400 $Y=1485 $D=89
M26 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6830 $Y=1485 $D=89
M27 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7260 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nand4_4 VNB VPB D C B A VPWR Y VGND
** N=92 EP=9 IP=0 FDC=32
*.SEEDPROM
M0 VGND D 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 10 D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND D 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 10 D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 11 C 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 10 C 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 11 C 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 10 C 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 11 B 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 12 B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 11 B 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5115 $Y=235 $D=9
M11 12 B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5535 $Y=235 $D=9
M12 Y A 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6015 $Y=235 $D=9
M13 12 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6435 $Y=235 $D=9
M14 Y A 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6855 $Y=235 $D=9
M15 12 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7275 $Y=235 $D=9
M16 Y D VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M17 VPWR D Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M18 Y D VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M19 VPWR D Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M20 Y C VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M21 VPWR C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M22 Y C VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M23 VPWR C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
M24 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4275 $Y=1485 $D=89
M25 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4695 $Y=1485 $D=89
M26 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5115 $Y=1485 $D=89
M27 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5535 $Y=1485 $D=89
M28 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6015 $Y=1485 $D=89
M29 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6435 $Y=1485 $D=89
M30 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6855 $Y=1485 $D=89
M31 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_4 VNB VPB A VPWR X VGND
** N=28 EP=6 IP=0 FDC=10
*.SEEDPROM
M0 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=885 $Y=235 $D=9
M2 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1315 $Y=235 $D=9
M3 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1745 $Y=235 $D=9
M4 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2175 $Y=235 $D=9
M5 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M6 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=880 $Y=1485 $D=89
M7 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1310 $Y=1485 $D=89
M8 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M9 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_1 VNB VPB A X VPWR VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND 7 X VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 7 A VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR 7 X VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 7 A VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__conb_1 HI VPWR VGND
** N=14 EP=3 IP=0 FDC=2
*.SEEDPROM
R0 HI VPWR 0.01 m=1 $[short] $X=105 $Y=1160 $D=284
R1 VGND LO 0.01 m=1 $[short] $X=795 $Y=1160 $D=284
.ENDS
***************************************
.SUBCKT ICV_90 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT CLK_RECOVERY VSS VDD CLK_OUT RESET_N BB_IN SCAN_IN<9> DATA_OUT SCAN_IN<10> SCAN_IN<21> SCAN_IN<20> SCAN_IN<8> SCAN_IN<18> SCAN_IN<7> CLK_IN SCAN_IN<19> SCAN_IN<11> SCAN_IN<12> SCAN_IN<15> SCAN_IN<14> SCAN_IN<16>
+ SCAN_IN<13> SCAN_IN<0> SCAN_IN<1> SCAN_IN<6> SCAN_IN<3> SCAN_IN<2> SCAN_IN<5> SCAN_IN<4> SCAN_IN<17>
** N=1147 EP=29 IP=15182 FDC=26384
M0 5 3 8 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=63950 $Y=84555 $D=9
M1 8 3 5 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=64370 $Y=84555 $D=9
M2 5 3 8 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=64790 $Y=84555 $D=9
M3 8 3 5 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=65210 $Y=84555 $D=9
M4 VSS CLK_OUT 8 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=65630 $Y=84555 $D=9
M5 8 CLK_OUT VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=66050 $Y=84555 $D=9
M6 VSS CLK_OUT 8 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=66470 $Y=84555 $D=9
M7 8 CLK_OUT VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=66890 $Y=84555 $D=9
M8 9 CLK_OUT VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=67840 $Y=84555 $D=9
M9 VSS CLK_OUT 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=68260 $Y=84555 $D=9
M10 9 CLK_OUT VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=68680 $Y=84555 $D=9
M11 VSS CLK_OUT 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=69100 $Y=84555 $D=9
M12 9 3 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=69520 $Y=84555 $D=9
M13 VSS 3 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=69940 $Y=84555 $D=9
M14 9 3 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=70360 $Y=84555 $D=9
M15 VSS 3 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=70780 $Y=84555 $D=9
M16 7 5 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=71740 $Y=84555 $D=9
M17 9 5 7 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=72160 $Y=84555 $D=9
M18 7 5 9 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=72580 $Y=84555 $D=9
M19 9 5 7 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=73000 $Y=84555 $D=9
M20 VDD 3 5 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=63950 $Y=85805 $D=89
M21 5 3 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=64370 $Y=85805 $D=89
M22 VDD 3 5 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=64790 $Y=85805 $D=89
M23 5 3 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=65210 $Y=85805 $D=89
M24 VDD CLK_OUT 5 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=65630 $Y=85805 $D=89
M25 5 CLK_OUT VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=66050 $Y=85805 $D=89
M26 VDD CLK_OUT 5 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=66470 $Y=85805 $D=89
M27 5 CLK_OUT VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=66890 $Y=85805 $D=89
M28 VDD CLK_OUT 6 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=67840 $Y=85805 $D=89
M29 6 CLK_OUT VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=68260 $Y=85805 $D=89
M30 VDD CLK_OUT 6 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=68680 $Y=85805 $D=89
M31 6 CLK_OUT VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=69100 $Y=85805 $D=89
M32 7 3 6 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=69520 $Y=85805 $D=89
M33 6 3 7 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=69940 $Y=85805 $D=89
M34 7 3 6 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=70360 $Y=85805 $D=89
M35 6 3 7 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=70780 $Y=85805 $D=89
M36 VDD 5 7 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=71740 $Y=85805 $D=89
M37 7 5 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=72160 $Y=85805 $D=89
M38 VDD 5 7 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=72580 $Y=85805 $D=89
M39 7 5 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=73000 $Y=85805 $D=89
X40 VSS VDD Dpar a=349.826 p=439.13 m=1 $[nwdiode] $X=5330 $Y=10690 $D=191
X41 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=14905 $D=191
X42 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=20345 $D=191
X43 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=25785 $D=191
X44 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=31225 $D=191
X45 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=36665 $D=191
X46 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=42105 $D=191
X47 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=47545 $D=191
X48 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=52985 $D=191
X49 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=58425 $D=191
X50 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=63865 $D=191
X51 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=69305 $D=191
X52 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=74745 $D=191
X53 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=80185 $D=191
X54 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=85625 $D=191
X55 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=91065 $D=191
X56 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=96505 $D=191
X57 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=101945 $D=191
X58 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=107385 $D=191
X59 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=112825 $D=191
X60 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=118265 $D=191
X61 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=123705 $D=191
X62 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=129145 $D=191
X63 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=134585 $D=191
X64 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=140025 $D=191
X65 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=145465 $D=191
X66 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=150905 $D=191
X67 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=156345 $D=191
X68 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=161785 $D=191
X69 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=167225 $D=191
X70 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=172665 $D=191
X71 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=178105 $D=191
X72 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=183545 $D=191
X73 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=188985 $D=191
X74 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=194425 $D=191
X75 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=199865 $D=191
X76 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=205305 $D=191
X77 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=210745 $D=191
X78 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=216185 $D=191
X79 VSS VDD Dpar a=616.827 p=441.58 m=1 $[nwdiode] $X=5330 $Y=221625 $D=191
X80 VSS VDD Dpar a=349.826 p=439.13 m=1 $[nwdiode] $X=5330 $Y=227065 $D=191
X81 1053 VDD Probe probetype=1 $[VDD] $X=114308 $Y=27288 $D=314
X82 1054 VSS Probe probetype=1 $[VSS] $X=114308 $Y=103878 $D=314
X83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 73440 1 0 $X=5330 $Y=70480
X84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 155040 0 0 $X=5330 $Y=154800
X85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 160480 0 0 $X=5330 $Y=160240
X86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 171360 1 0 $X=5330 $Y=168400
X87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 198560 1 0 $X=5330 $Y=195600
X88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 225760 0 0 $X=5330 $Y=225520
X89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=6900 133280 1 0 $X=6710 $Y=130320
X90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=9200 149600 0 0 $X=9010 $Y=149360
X91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=19320 13600 0 0 $X=19130 $Y=13360
X92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=25300 127840 1 0 $X=25110 $Y=124880
X93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=25760 68000 1 0 $X=25570 $Y=65040
X94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=31280 144160 1 0 $X=31090 $Y=141200
X95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=32200 29920 1 0 $X=32010 $Y=26960
X96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=34040 19040 0 0 $X=33850 $Y=18800
X97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=34040 46240 0 0 $X=33850 $Y=46000
X98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=34960 106080 1 0 $X=34770 $Y=103120
X99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=35420 78880 1 0 $X=35230 $Y=75920
X100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=38640 62560 1 0 $X=38450 $Y=59600
X101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=48300 73440 1 0 $X=48110 $Y=70480
X102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=48300 111520 1 0 $X=48110 $Y=108560
X103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=51060 209440 1 0 $X=50870 $Y=206480
X104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=52900 198560 0 0 $X=52710 $Y=198320
X105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=55660 29920 1 0 $X=55470 $Y=26960
X106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=55660 127840 1 0 $X=55470 $Y=124880
X107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=62100 84320 0 0 $X=61910 $Y=84080
X108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=74980 122400 0 0 $X=74790 $Y=122160
X109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=83260 51680 1 0 $X=83070 $Y=48720
X110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=86940 149600 1 0 $X=86750 $Y=146640
X111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=104420 89760 1 0 $X=104230 $Y=86800
X112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=104880 78880 0 0 $X=104690 $Y=78640
X113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=108560 89760 0 0 $X=108370 $Y=89520
X114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=117760 84320 1 0 $X=117570 $Y=81360
X115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=122360 116960 1 0 $X=122170 $Y=114000
X116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=127420 198560 1 0 $X=127230 $Y=195600
X117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=129260 100640 0 0 $X=129070 $Y=100400
X118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=136160 155040 0 0 $X=135970 $Y=154800
X119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=143060 171360 1 0 $X=142870 $Y=168400
X120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=146280 160480 0 0 $X=146090 $Y=160240
X121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=147200 127840 1 0 $X=147010 $Y=124880
X122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=160540 35360 1 0 $X=160350 $Y=32400
X123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=160540 62560 1 0 $X=160350 $Y=59600
X124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=163760 133280 0 0 $X=163570 $Y=133040
X125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=172960 24480 1 0 $X=172770 $Y=21520
X126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=175720 127840 1 0 $X=175530 $Y=124880
X127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=188600 187680 1 0 $X=188410 $Y=184720
X128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=189520 193120 0 0 $X=189330 $Y=192880
X129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=191360 165920 1 0 $X=191170 $Y=162960
X130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=194120 24480 1 0 $X=193930 $Y=21520
X131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=194120 111520 1 0 $X=193930 $Y=108560
X132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=194120 220320 1 0 $X=193930 $Y=217360
X133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=198260 209440 1 0 $X=198070 $Y=206480
X134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=198720 95200 1 0 $X=198530 $Y=92240
X135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=200560 176800 0 0 $X=200370 $Y=176560
X136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=202400 73440 0 0 $X=202210 $Y=73200
X137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=203320 198560 1 0 $X=203130 $Y=195600
X138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=205160 193120 1 0 $X=204970 $Y=190160
X139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=220340 133280 0 0 $X=220150 $Y=133040
X140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 13600 0 180 $X=221530 $Y=10640
X141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 29920 0 180 $X=221530 $Y=26960
X142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 57120 0 180 $X=221530 $Y=54160
X143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 62560 0 180 $X=221530 $Y=59600
X144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 89760 0 180 $X=221530 $Y=86800
X145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 116960 0 180 $X=221530 $Y=114000
X146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 127840 0 180 $X=221530 $Y=124880
X147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 155040 0 180 $X=221530 $Y=152080
X148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 160480 0 180 $X=221530 $Y=157520
X149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 165920 0 180 $X=221530 $Y=162960
X150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 171360 0 180 $X=221530 $Y=168400
X151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 187680 0 180 $X=221530 $Y=184720
X152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 198560 0 180 $X=221530 $Y=195600
X153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 209440 0 180 $X=221530 $Y=206480
X154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=223100 225760 1 180 $X=221530 $Y=225520
X155 VSS VDD ICV_1 $T=5520 62560 0 0 $X=5330 $Y=62320
X156 VSS VDD ICV_1 $T=5520 149600 0 0 $X=5330 $Y=149360
X157 VSS VDD ICV_1 $T=6900 51680 0 0 $X=6710 $Y=51440
X158 VSS VDD ICV_1 $T=6900 84320 0 0 $X=6710 $Y=84080
X159 VSS VDD ICV_1 $T=223100 116960 1 180 $X=221530 $Y=116720
X160 VSS VDD ICV_1 $T=223100 187680 1 180 $X=221530 $Y=187440
X161 VSS VDD ICV_1 $T=223100 198560 1 180 $X=221530 $Y=198320
X162 VSS VDD ICV_1 $T=223100 220320 1 180 $X=221530 $Y=220080
X163 VSS VDD ICV_2 $T=5520 138720 0 0 $X=5330 $Y=138480
X164 VSS VDD ICV_2 $T=223100 13600 1 180 $X=221530 $Y=13360
X165 VSS VDD ICV_2 $T=223100 171360 1 180 $X=221530 $Y=171120
X166 VSS VDD ICV_2 $T=223100 209440 1 180 $X=221530 $Y=209200
X167 VSS VDD ICV_3 $T=5520 19040 0 0 $X=5330 $Y=18800
X168 VSS VDD ICV_3 $T=5520 40800 0 0 $X=5330 $Y=40560
X169 VSS VDD ICV_3 $T=5520 73440 0 0 $X=5330 $Y=73200
X170 VSS VDD ICV_3 $T=5520 95200 0 0 $X=5330 $Y=94960
X171 VSS VDD ICV_3 $T=5520 116960 0 0 $X=5330 $Y=116720
X172 VSS VDD ICV_3 $T=5520 171360 0 0 $X=5330 $Y=171120
X173 VSS VDD ICV_3 $T=5520 198560 0 0 $X=5330 $Y=198320
X174 VSS VDD ICV_3 $T=223100 29920 1 180 $X=221530 $Y=29680
X175 VSS VDD ICV_3 $T=223100 62560 1 180 $X=221530 $Y=62320
X176 VSS VDD ICV_3 $T=223100 89760 1 180 $X=221530 $Y=89520
X177 VSS VDD ICV_3 $T=223100 127840 1 180 $X=221530 $Y=127600
X250 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=21620 193120 0 0 $X=21430 $Y=192880
X251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=27600 73440 1 0 $X=27410 $Y=70480
X252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=28520 149600 0 0 $X=28330 $Y=149360
X253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=29440 19040 0 0 $X=29250 $Y=18800
X254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=37720 193120 1 0 $X=37530 $Y=190160
X255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=40020 73440 1 0 $X=39830 $Y=70480
X256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=41400 106080 0 0 $X=41210 $Y=105840
X257 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=47380 106080 0 0 $X=47190 $Y=105840
X258 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=48300 40800 1 0 $X=48110 $Y=37840
X259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=48300 155040 1 0 $X=48110 $Y=152080
X260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=54740 78880 0 0 $X=54550 $Y=78640
X261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=59800 176800 1 0 $X=59610 $Y=173840
X262 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=60720 111520 1 0 $X=60530 $Y=108560
X263 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=61180 133280 1 0 $X=60990 $Y=130320
X264 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=76360 40800 1 0 $X=76170 $Y=37840
X265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=81420 111520 0 0 $X=81230 $Y=111280
X266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=83720 187680 1 0 $X=83530 $Y=184720
X267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=85560 160480 0 0 $X=85370 $Y=160240
X268 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=87400 160480 1 0 $X=87210 $Y=157520
X269 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=102120 95200 0 0 $X=101930 $Y=94960
X270 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=103040 127840 0 0 $X=102850 $Y=127600
X271 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=104420 84320 1 0 $X=104230 $Y=81360
X272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=113620 35360 0 0 $X=113430 $Y=35120
X273 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=115920 160480 1 0 $X=115730 $Y=157520
X274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=121440 111520 1 0 $X=121250 $Y=108560
X275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=126040 78880 1 0 $X=125850 $Y=75920
X276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=139840 35360 0 0 $X=139650 $Y=35120
X277 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=139840 220320 0 0 $X=139650 $Y=220080
X278 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=140760 78880 0 0 $X=140570 $Y=78640
X279 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=155940 84320 1 0 $X=155750 $Y=81360
X280 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=157780 40800 1 0 $X=157590 $Y=37840
X281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=158700 84320 0 0 $X=158510 $Y=84080
X282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=163300 116960 0 0 $X=163110 $Y=116720
X283 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=166980 57120 0 0 $X=166790 $Y=56880
X284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=169740 182240 0 0 $X=169550 $Y=182000
X285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=169740 220320 0 0 $X=169550 $Y=220080
X286 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=174340 78880 1 0 $X=174150 $Y=75920
X287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=174340 214880 0 0 $X=174150 $Y=214640
X288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=176640 57120 1 0 $X=176450 $Y=54160
X289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=181240 144160 1 0 $X=181050 $Y=141200
X290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=182620 149600 1 0 $X=182430 $Y=146640
X291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=183540 19040 1 0 $X=183350 $Y=16080
X292 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=188600 127840 1 0 $X=188410 $Y=124880
X293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=188600 133280 1 0 $X=188410 $Y=130320
X294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=199180 106080 1 0 $X=198990 $Y=103120
X295 VSS VDD ICV_4 $T=19780 182240 1 0 $X=19590 $Y=179280
X296 VSS VDD ICV_4 $T=19780 187680 1 0 $X=19590 $Y=184720
X297 VSS VDD ICV_4 $T=33580 198560 0 0 $X=33390 $Y=198320
X298 VSS VDD ICV_4 $T=47840 220320 1 0 $X=47650 $Y=217360
X299 VSS VDD ICV_4 $T=75900 62560 1 0 $X=75710 $Y=59600
X300 VSS VDD ICV_4 $T=75900 138720 1 0 $X=75710 $Y=135760
X301 VSS VDD ICV_4 $T=89700 95200 0 0 $X=89510 $Y=94960
X302 VSS VDD ICV_4 $T=89700 106080 0 0 $X=89510 $Y=105840
X303 VSS VDD ICV_4 $T=89700 133280 0 0 $X=89510 $Y=133040
X304 VSS VDD ICV_4 $T=89700 138720 0 0 $X=89510 $Y=138480
X305 VSS VDD ICV_4 $T=89700 144160 0 0 $X=89510 $Y=143920
X306 VSS VDD ICV_4 $T=103960 220320 1 0 $X=103770 $Y=217360
X307 VSS VDD ICV_4 $T=117760 68000 0 0 $X=117570 $Y=67760
X308 VSS VDD ICV_4 $T=117760 176800 0 0 $X=117570 $Y=176560
X309 VSS VDD ICV_4 $T=145820 193120 0 0 $X=145630 $Y=192880
X310 VSS VDD ICV_4 $T=160080 40800 1 0 $X=159890 $Y=37840
X311 VSS VDD ICV_4 $T=160080 133280 1 0 $X=159890 $Y=130320
X312 VSS VDD ICV_4 $T=173880 51680 0 0 $X=173690 $Y=51440
X313 VSS VDD ICV_4 $T=173880 62560 0 0 $X=173690 $Y=62320
X314 VSS VDD ICV_4 $T=173880 193120 0 0 $X=173690 $Y=192880
X315 VSS VDD ICV_4 $T=188140 68000 1 0 $X=187950 $Y=65040
X316 VSS VDD ICV_4 $T=188140 78880 1 0 $X=187950 $Y=75920
X317 VSS VDD ICV_4 $T=188140 204000 1 0 $X=187950 $Y=201040
X318 VSS VDD ICV_4 $T=201940 68000 0 0 $X=201750 $Y=67760
X319 VSS VDD ICV_4 $T=201940 220320 0 0 $X=201750 $Y=220080
X320 VSS VDD ICV_4 $T=219420 13600 1 0 $X=219230 $Y=10640
X321 VSS VDD ICV_4 $T=219420 225760 0 0 $X=219230 $Y=225520
X322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 40800 1 0 $X=6710 $Y=37840
X323 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 57120 0 0 $X=6710 $Y=56880
X324 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 198560 0 0 $X=6710 $Y=198320
X325 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=16560 187680 1 0 $X=16370 $Y=184720
X326 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=18400 122400 0 0 $X=18210 $Y=122160
X327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=20240 73440 1 0 $X=20050 $Y=70480
X328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=25760 62560 1 0 $X=25570 $Y=59600
X329 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=27600 40800 1 0 $X=27410 $Y=37840
X330 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=28060 165920 1 0 $X=27870 $Y=162960
X331 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=28060 193120 1 0 $X=27870 $Y=190160
X332 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=31280 13600 1 0 $X=31090 $Y=10640
X333 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=34040 73440 0 0 $X=33850 $Y=73200
X334 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=36340 84320 1 0 $X=36150 $Y=81360
X335 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=50600 116960 0 0 $X=50410 $Y=116720
X336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=58420 138720 0 0 $X=58230 $Y=138480
X337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=62100 106080 0 0 $X=61910 $Y=105840
X338 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=63020 95200 1 0 $X=62830 $Y=92240
X339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=63020 100640 1 0 $X=62830 $Y=97680
X340 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=65780 40800 0 0 $X=65590 $Y=40560
X341 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=65780 57120 1 0 $X=65590 $Y=54160
X342 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=66700 182240 1 0 $X=66510 $Y=179280
X343 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=68540 198560 0 0 $X=68350 $Y=198320
X344 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=76360 106080 1 0 $X=76170 $Y=103120
X345 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=78200 182240 1 0 $X=78010 $Y=179280
X346 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=81420 95200 1 0 $X=81230 $Y=92240
X347 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=82800 193120 1 0 $X=82610 $Y=190160
X348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=83720 24480 1 0 $X=83530 $Y=21520
X349 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=85100 100640 0 0 $X=84910 $Y=100400
X350 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=85100 144160 1 0 $X=84910 $Y=141200
X351 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=86940 182240 1 0 $X=86750 $Y=179280
X352 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=90160 68000 0 0 $X=89970 $Y=67760
X353 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=90620 68000 1 0 $X=90430 $Y=65040
X354 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=92000 209440 0 0 $X=91810 $Y=209200
X355 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=95680 46240 1 0 $X=95490 $Y=43280
X356 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=96600 35360 1 0 $X=96410 $Y=32400
X357 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=98440 24480 1 0 $X=98250 $Y=21520
X358 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=99360 176800 1 0 $X=99170 $Y=173840
X359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=101660 155040 0 0 $X=101470 $Y=154800
X360 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=104420 40800 1 0 $X=104230 $Y=37840
X361 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=108560 214880 1 0 $X=108370 $Y=211920
X362 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=114540 68000 0 0 $X=114350 $Y=67760
X363 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=114540 73440 0 0 $X=114350 $Y=73200
X364 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=115460 155040 1 0 $X=115270 $Y=152080
X365 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=121900 149600 0 0 $X=121710 $Y=149360
X366 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=129260 51680 0 0 $X=129070 $Y=51440
X367 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=129260 111520 0 0 $X=129070 $Y=111280
X368 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=134320 68000 1 0 $X=134130 $Y=65040
X369 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=134320 160480 1 0 $X=134130 $Y=157520
X370 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=136620 193120 1 0 $X=136430 $Y=190160
X371 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=137540 57120 1 0 $X=137350 $Y=54160
X372 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=139840 144160 1 0 $X=139650 $Y=141200
X373 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=140760 220320 1 0 $X=140570 $Y=217360
X374 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=141220 51680 0 0 $X=141030 $Y=51440
X375 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=141680 160480 1 0 $X=141490 $Y=157520
X376 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=147660 51680 1 0 $X=147470 $Y=48720
X377 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=151340 78880 1 0 $X=151150 $Y=75920
X378 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=151800 84320 1 0 $X=151610 $Y=81360
X379 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=151800 111520 0 0 $X=151610 $Y=111280
X380 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=153640 95200 0 0 $X=153450 $Y=94960
X381 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=156860 193120 1 0 $X=156670 $Y=190160
X382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=164680 19040 1 0 $X=164490 $Y=16080
X383 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=166060 122400 1 0 $X=165870 $Y=119440
X384 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=171120 171360 0 0 $X=170930 $Y=171120
X385 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=178480 84320 0 0 $X=178290 $Y=84080
X386 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=188140 225760 0 0 $X=187950 $Y=225520
X387 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=190440 225760 1 0 $X=190250 $Y=222800
X388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=190900 149600 1 0 $X=190710 $Y=146640
X389 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=191360 176800 0 0 $X=191170 $Y=176560
X390 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=192740 100640 1 0 $X=192550 $Y=97680
X391 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=192740 198560 1 0 $X=192550 $Y=195600
X392 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=195040 106080 1 0 $X=194850 $Y=103120
X393 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=195500 35360 1 0 $X=195310 $Y=32400
X394 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=195960 138720 1 0 $X=195770 $Y=135760
X395 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=216660 225760 0 0 $X=216470 $Y=225520
X396 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=218960 204000 1 0 $X=218770 $Y=201040
X397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=6900 176800 0 0 $X=6710 $Y=176560
X398 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=13800 198560 1 0 $X=13610 $Y=195600
X399 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=15640 78880 1 0 $X=15450 $Y=75920
X400 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=18400 144160 0 0 $X=18210 $Y=143920
X401 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=27600 176800 0 0 $X=27410 $Y=176560
X402 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=28060 138720 0 0 $X=27870 $Y=138480
X403 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=29900 35360 1 0 $X=29710 $Y=32400
X404 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=34040 51680 0 0 $X=33850 $Y=51440
X405 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=40480 160480 1 0 $X=40290 $Y=157520
X406 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=40940 171360 1 0 $X=40750 $Y=168400
X407 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43240 89760 1 0 $X=43050 $Y=86800
X408 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43700 138720 0 0 $X=43510 $Y=138480
X409 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43700 225760 1 0 $X=43510 $Y=222800
X410 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=47380 204000 0 0 $X=47190 $Y=203760
X411 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=48300 29920 1 0 $X=48110 $Y=26960
X412 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=50600 204000 1 0 $X=50410 $Y=201040
X413 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=55660 209440 0 0 $X=55470 $Y=209200
X414 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=59340 116960 1 0 $X=59150 $Y=114000
X415 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=63480 193120 1 0 $X=63290 $Y=190160
X416 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=64860 46240 1 0 $X=64670 $Y=43280
X417 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=69460 155040 1 0 $X=69270 $Y=152080
X418 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=72220 220320 1 0 $X=72030 $Y=217360
X419 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=74980 57120 0 0 $X=74790 $Y=56880
X420 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=75440 62560 0 0 $X=75250 $Y=62320
X421 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=78660 19040 1 0 $X=78470 $Y=16080
X422 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=79120 51680 0 0 $X=78930 $Y=51440
X423 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=80500 57120 1 0 $X=80310 $Y=54160
X424 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=80500 84320 1 0 $X=80310 $Y=81360
X425 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=82800 19040 0 0 $X=82610 $Y=18800
X426 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=82800 214880 1 0 $X=82610 $Y=211920
X427 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=85100 29920 0 0 $X=84910 $Y=29680
X428 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=91540 100640 1 0 $X=91350 $Y=97680
X429 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=92460 209440 1 0 $X=92270 $Y=206480
X430 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=93840 35360 0 0 $X=93650 $Y=35120
X431 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=96600 144160 1 0 $X=96410 $Y=141200
X432 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=97060 204000 1 0 $X=96870 $Y=201040
X433 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=100280 116960 0 0 $X=100090 $Y=116720
X434 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=107640 24480 0 0 $X=107450 $Y=24240
X435 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=110400 116960 0 0 $X=110210 $Y=116720
X436 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=112700 225760 1 0 $X=112510 $Y=222800
X437 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=114080 220320 1 0 $X=113890 $Y=217360
X438 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=114540 116960 1 0 $X=114350 $Y=114000
X439 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=119140 106080 1 0 $X=118950 $Y=103120
X440 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=121440 35360 1 0 $X=121250 $Y=32400
X441 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=123280 122400 1 0 $X=123090 $Y=119440
X442 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=129260 204000 0 0 $X=129070 $Y=203760
X443 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=132480 127840 1 0 $X=132290 $Y=124880
X444 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=132940 62560 0 0 $X=132750 $Y=62320
X445 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=132940 116960 0 0 $X=132750 $Y=116720
X446 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=134780 95200 1 0 $X=134590 $Y=92240
X447 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=139380 46240 1 0 $X=139190 $Y=43280
X448 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=142600 133280 1 0 $X=142410 $Y=130320
X449 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=148120 214880 1 0 $X=147930 $Y=211920
X450 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=148580 149600 1 0 $X=148390 $Y=146640
X451 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=152260 144160 1 0 $X=152070 $Y=141200
X452 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=153180 176800 1 0 $X=152990 $Y=173840
X453 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=153640 19040 1 0 $X=153450 $Y=16080
X454 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=154100 122400 1 0 $X=153910 $Y=119440
X455 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=155940 187680 1 0 $X=155750 $Y=184720
X456 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=163300 122400 0 0 $X=163110 $Y=122160
X457 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=163760 209440 0 0 $X=163570 $Y=209200
X458 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=164680 214880 0 0 $X=164490 $Y=214640
X459 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=166060 84320 0 0 $X=165870 $Y=84080
X460 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=166520 46240 0 0 $X=166330 $Y=46000
X461 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=167440 84320 1 0 $X=167250 $Y=81360
X462 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=168360 149600 1 0 $X=168170 $Y=146640
X463 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=172040 68000 1 0 $X=171850 $Y=65040
X464 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=172500 29920 1 0 $X=172310 $Y=26960
X465 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=173880 73440 1 0 $X=173690 $Y=70480
X466 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=174340 19040 1 0 $X=174150 $Y=16080
X467 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=184460 78880 1 0 $X=184270 $Y=75920
X468 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=195960 165920 1 0 $X=195770 $Y=162960
X469 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=196420 68000 1 0 $X=196230 $Y=65040
X470 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=197340 24480 0 0 $X=197150 $Y=24240
X471 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=201940 116960 1 0 $X=201750 $Y=114000
X472 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=202400 122400 1 0 $X=202210 $Y=119440
X473 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=202400 144160 1 0 $X=202210 $Y=141200
X474 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=202400 182240 1 0 $X=202210 $Y=179280
X475 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=207000 209440 1 0 $X=206810 $Y=206480
X476 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=217120 40800 0 0 $X=216930 $Y=40560
X477 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=217120 62560 0 0 $X=216930 $Y=62320
X478 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=217120 209440 0 0 $X=216930 $Y=209200
X479 VSS VDD ICV_5 $T=218040 24480 0 0 $X=217850 $Y=24240
X480 VSS VDD ICV_5 $T=218040 51680 0 0 $X=217850 $Y=51440
X481 VSS VDD ICV_5 $T=218040 57120 0 0 $X=217850 $Y=56880
X482 VSS VDD ICV_5 $T=218040 84320 0 0 $X=217850 $Y=84080
X483 VSS VDD ICV_5 $T=218040 111520 0 0 $X=217850 $Y=111280
X484 VSS VDD ICV_5 $T=218040 122400 0 0 $X=217850 $Y=122160
X485 VSS VDD ICV_5 $T=218040 149600 0 0 $X=217850 $Y=149360
X486 VSS VDD ICV_5 $T=218040 155040 0 0 $X=217850 $Y=154800
X487 VSS VDD ICV_5 $T=218040 160480 0 0 $X=217850 $Y=160240
X488 VSS VDD ICV_5 $T=218040 165920 0 0 $X=217850 $Y=165680
X489 VSS VDD ICV_5 $T=218040 182240 0 0 $X=217850 $Y=182000
X490 VSS VDD ICV_5 $T=218040 193120 0 0 $X=217850 $Y=192880
X491 VSS VDD ICV_5 $T=218040 204000 0 0 $X=217850 $Y=203760
X492 VSS VDD 62 VDD 61 VSS sky130_fd_sc_hd__buf_1 $T=12420 35360 0 0 $X=12230 $Y=35120
X493 VSS VDD 57 VDD 87 VSS sky130_fd_sc_hd__buf_1 $T=13800 176800 0 0 $X=13610 $Y=176560
X494 VSS VDD 108 VDD 24 VSS sky130_fd_sc_hd__buf_1 $T=18860 62560 0 0 $X=18670 $Y=62320
X495 VSS VDD 120 VDD 26 VSS sky130_fd_sc_hd__buf_1 $T=26680 95200 0 0 $X=26490 $Y=94960
X496 VSS VDD 164 VDD 43 VSS sky130_fd_sc_hd__buf_1 $T=27140 68000 0 0 $X=26950 $Y=67760
X497 VSS VDD 148 VDD 173 VSS sky130_fd_sc_hd__buf_1 $T=28060 160480 1 0 $X=27870 $Y=157520
X498 VSS VDD 153 VDD 119 VSS sky130_fd_sc_hd__buf_1 $T=28980 62560 1 0 $X=28790 $Y=59600
X499 VSS VDD 204 VDD 210 VSS sky130_fd_sc_hd__buf_1 $T=34960 62560 1 0 $X=34770 $Y=59600
X500 VSS VDD 184 VDD 58 VSS sky130_fd_sc_hd__buf_1 $T=34960 204000 0 0 $X=34770 $Y=203760
X501 VSS VDD 184 VDD 166 VSS sky130_fd_sc_hd__buf_1 $T=36340 220320 1 0 $X=36150 $Y=217360
X502 VSS VDD 161 VDD 190 VSS sky130_fd_sc_hd__buf_1 $T=37260 187680 0 0 $X=37070 $Y=187440
X503 VSS VDD 225 VDD 106 VSS sky130_fd_sc_hd__buf_1 $T=39100 209440 1 0 $X=38910 $Y=206480
X504 VSS VDD 230 VDD 187 VSS sky130_fd_sc_hd__buf_1 $T=39560 144160 0 0 $X=39370 $Y=143920
X505 VSS VDD 206 VDD 189 VSS sky130_fd_sc_hd__buf_1 $T=39560 193120 1 0 $X=39370 $Y=190160
X506 VSS VDD 188 VDD 231 VSS sky130_fd_sc_hd__buf_1 $T=42780 144160 1 0 $X=42590 $Y=141200
X507 VSS VDD 206 VDD 240 VSS sky130_fd_sc_hd__buf_1 $T=42780 198560 0 0 $X=42590 $Y=198320
X508 VSS VDD 259 VDD 232 VSS sky130_fd_sc_hd__buf_1 $T=49220 24480 1 0 $X=49030 $Y=21520
X509 VSS VDD 248 VDD 109 VSS sky130_fd_sc_hd__buf_1 $T=49220 149600 1 0 $X=49030 $Y=146640
X510 VSS VDD 249 VDD 271 VSS sky130_fd_sc_hd__buf_1 $T=49220 187680 1 0 $X=49030 $Y=184720
X511 VSS VDD 302 VDD 250 VSS sky130_fd_sc_hd__buf_1 $T=52440 35360 1 0 $X=52250 $Y=32400
X512 VSS VDD 17 VDD 281 VSS sky130_fd_sc_hd__buf_1 $T=53360 111520 0 0 $X=53170 $Y=111280
X513 VSS VDD 301 VDD 145 VSS sky130_fd_sc_hd__buf_1 $T=60260 214880 1 0 $X=60070 $Y=211920
X514 VSS VDD 272 VDD 357 VSS sky130_fd_sc_hd__buf_1 $T=63020 209440 0 0 $X=62830 $Y=209200
X515 VSS VDD 324 VDD 339 VSS sky130_fd_sc_hd__buf_1 $T=63480 171360 1 0 $X=63290 $Y=168400
X516 VSS VDD 372 VDD 128 VSS sky130_fd_sc_hd__buf_1 $T=67620 40800 1 0 $X=67430 $Y=37840
X517 VSS VDD 355 VDD 188 VSS sky130_fd_sc_hd__buf_1 $T=68080 133280 1 0 $X=67890 $Y=130320
X518 VSS VDD 382 VDD 317 VSS sky130_fd_sc_hd__buf_1 $T=69920 19040 1 0 $X=69730 $Y=16080
X519 VSS VDD 150 VDD 401 VSS sky130_fd_sc_hd__buf_1 $T=71760 198560 0 0 $X=71570 $Y=198320
X520 VSS VDD 400 VDD 348 VSS sky130_fd_sc_hd__buf_1 $T=74060 149600 0 0 $X=73870 $Y=149360
X521 VSS VDD 388 VDD 356 VSS sky130_fd_sc_hd__buf_1 $T=76360 122400 0 0 $X=76170 $Y=122160
X522 VSS VDD 326 VDD 158 VSS sky130_fd_sc_hd__buf_1 $T=84640 106080 0 0 $X=84450 $Y=105840
X523 VSS VDD 326 VDD 466 VSS sky130_fd_sc_hd__buf_1 $T=91080 100640 0 0 $X=90890 $Y=100400
X524 VSS VDD 17 VDD 473 VSS sky130_fd_sc_hd__buf_1 $T=91540 89760 0 0 $X=91350 $Y=89520
X525 VSS VDD 17 VDD 346 VSS sky130_fd_sc_hd__buf_1 $T=92000 106080 1 0 $X=91810 $Y=103120
X526 VSS VDD 377 VDD 337 VSS sky130_fd_sc_hd__buf_1 $T=92000 160480 0 0 $X=91810 $Y=160240
X527 VSS VDD 505 VDD 492 VSS sky130_fd_sc_hd__buf_1 $T=96600 225760 1 0 $X=96410 $Y=222800
X528 VSS VDD 509 VDD 393 VSS sky130_fd_sc_hd__buf_1 $T=98900 89760 1 0 $X=98710 $Y=86800
X529 VSS VDD 509 VDD 458 VSS sky130_fd_sc_hd__buf_1 $T=104420 84320 0 0 $X=104230 $Y=84080
X530 VSS VDD 522 VDD 489 VSS sky130_fd_sc_hd__buf_1 $T=109940 35360 1 0 $X=109750 $Y=32400
X531 VSS VDD 554 VDD 522 VSS sky130_fd_sc_hd__buf_1 $T=111780 19040 0 0 $X=111590 $Y=18800
X532 VSS VDD 534 VDD 529 VSS sky130_fd_sc_hd__buf_1 $T=111780 57120 0 0 $X=111590 $Y=56880
X533 VSS VDD 573 VDD 565 VSS sky130_fd_sc_hd__buf_1 $T=112700 84320 0 0 $X=112510 $Y=84080
X534 VSS VDD 604 VDD 534 VSS sky130_fd_sc_hd__buf_1 $T=115460 51680 1 0 $X=115270 $Y=48720
X535 VSS VDD 630 VDD 605 VSS sky130_fd_sc_hd__buf_1 $T=119140 138720 1 0 $X=118950 $Y=135760
X536 VSS VDD 600 VDD 635 VSS sky130_fd_sc_hd__buf_1 $T=119140 171360 1 0 $X=118950 $Y=168400
X537 VSS VDD 632 VDD 623 VSS sky130_fd_sc_hd__buf_1 $T=131560 40800 0 0 $X=131370 $Y=40560
X538 VSS VDD 666 VDD 628 VSS sky130_fd_sc_hd__buf_1 $T=133400 24480 1 0 $X=133210 $Y=21520
X539 VSS VDD 673 VDD 620 VSS sky130_fd_sc_hd__buf_1 $T=136620 165920 0 0 $X=136430 $Y=165680
X540 VSS VDD 622 VDD 703 VSS sky130_fd_sc_hd__buf_1 $T=140300 57120 1 0 $X=140110 $Y=54160
X541 VSS VDD 578 VDD 730 VSS sky130_fd_sc_hd__buf_1 $T=140300 62560 1 0 $X=140110 $Y=59600
X542 VSS VDD 700 VDD 676 VSS sky130_fd_sc_hd__buf_1 $T=140760 19040 0 0 $X=140570 $Y=18800
X543 VSS VDD 719 VDD 519 VSS sky130_fd_sc_hd__buf_1 $T=140760 29920 0 0 $X=140570 $Y=29680
X544 VSS VDD 509 VDD 701 VSS sky130_fd_sc_hd__buf_1 $T=140760 73440 0 0 $X=140570 $Y=73200
X545 VSS VDD 752 VDD 641 VSS sky130_fd_sc_hd__buf_1 $T=146280 204000 1 0 $X=146090 $Y=201040
X546 VSS VDD 744 VDD 574 VSS sky130_fd_sc_hd__buf_1 $T=147200 46240 0 0 $X=147010 $Y=46000
X547 VSS VDD 731 VDD 783 VSS sky130_fd_sc_hd__buf_1 $T=149960 78880 1 0 $X=149770 $Y=75920
X548 VSS VDD 770 VDD 471 VSS sky130_fd_sc_hd__buf_1 $T=151340 204000 1 0 $X=151150 $Y=201040
X549 VSS VDD 789 VDD 674 VSS sky130_fd_sc_hd__buf_1 $T=152260 29920 1 0 $X=152070 $Y=26960
X550 VSS VDD 677 VDD 596 VSS sky130_fd_sc_hd__buf_1 $T=152720 73440 0 0 $X=152530 $Y=73200
X551 VSS VDD 520 VDD 787 VSS sky130_fd_sc_hd__buf_1 $T=153640 78880 0 0 $X=153450 $Y=78640
X552 VSS VDD 783 VDD 698 VSS sky130_fd_sc_hd__buf_1 $T=154560 84320 1 0 $X=154370 $Y=81360
X553 VSS VDD 677 VDD 521 VSS sky130_fd_sc_hd__buf_1 $T=155020 116960 1 0 $X=154830 $Y=114000
X554 VSS VDD 798 VDD 537 VSS sky130_fd_sc_hd__buf_1 $T=156860 193120 0 0 $X=156670 $Y=192880
X555 VSS VDD 823 VDD 690 VSS sky130_fd_sc_hd__buf_1 $T=161460 209440 1 0 $X=161270 $Y=206480
X556 VSS VDD 846 VDD 745 VSS sky130_fd_sc_hd__buf_1 $T=165140 138720 1 0 $X=164950 $Y=135760
X557 VSS VDD 865 VDD 788 VSS sky130_fd_sc_hd__buf_1 $T=168820 24480 0 0 $X=168630 $Y=24240
X558 VSS VDD 872 VDD 819 VSS sky130_fd_sc_hd__buf_1 $T=171120 171360 1 0 $X=170930 $Y=168400
X559 VSS VDD 878 VDD 865 VSS sky130_fd_sc_hd__buf_1 $T=171580 24480 1 0 $X=171390 $Y=21520
X560 VSS VDD 765 VDD 756 VSS sky130_fd_sc_hd__buf_1 $T=176180 68000 1 0 $X=175990 $Y=65040
X561 VSS VDD 749 VDD 902 VSS sky130_fd_sc_hd__buf_1 $T=181240 57120 1 0 $X=181050 $Y=54160
X562 VSS VDD 910 VDD 769 VSS sky130_fd_sc_hd__buf_1 $T=181240 149600 1 0 $X=181050 $Y=146640
X563 VSS VDD 904 VDD 830 VSS sky130_fd_sc_hd__buf_1 $T=182620 24480 1 0 $X=182430 $Y=21520
X564 VSS VDD 946 VDD 547 VSS sky130_fd_sc_hd__buf_1 $T=188140 187680 0 0 $X=187950 $Y=187440
X565 VSS VDD 947 VDD 913 VSS sky130_fd_sc_hd__buf_1 $T=190900 193120 0 0 $X=190710 $Y=192880
X566 VSS VDD 967 VDD 892 VSS sky130_fd_sc_hd__buf_1 $T=193660 127840 1 0 $X=193470 $Y=124880
X567 VSS VDD 956 VDD 912 VSS sky130_fd_sc_hd__buf_1 $T=194120 73440 0 0 $X=193930 $Y=73200
X568 VSS VDD 935 VDD 760 VSS sky130_fd_sc_hd__buf_1 $T=196420 29920 0 0 $X=196230 $Y=29680
X569 VSS VDD 650 VDD 985 VSS sky130_fd_sc_hd__buf_1 $T=196880 68000 0 0 $X=196690 $Y=67760
X570 VSS VDD 960 VDD 928 VSS sky130_fd_sc_hd__buf_1 $T=196880 155040 0 0 $X=196690 $Y=154800
X571 VSS VDD 987 VDD 774 VSS sky130_fd_sc_hd__buf_1 $T=197800 106080 1 0 $X=197610 $Y=103120
X572 VSS VDD 940 VDD 721 VSS sky130_fd_sc_hd__buf_1 $T=198720 138720 1 0 $X=198530 $Y=135760
X573 VSS VDD 1003 VDD 757 VSS sky130_fd_sc_hd__buf_1 $T=200560 127840 1 0 $X=200370 $Y=124880
X574 VSS VDD 972 VDD 988 VSS sky130_fd_sc_hd__buf_1 $T=203320 122400 0 0 $X=203130 $Y=122160
X575 VSS VDD 1019 VDD 914 VSS sky130_fd_sc_hd__buf_1 $T=207000 100640 0 0 $X=206810 $Y=100400
X576 VSS VDD 1034 VDD 963 VSS sky130_fd_sc_hd__buf_1 $T=211140 73440 1 0 $X=210950 $Y=70480
X577 VSS VDD 1033 VDD 851 VSS sky130_fd_sc_hd__buf_1 $T=217580 204000 1 0 $X=217390 $Y=201040
X578 VSS 20 sky130_fd_sc_hd__diode_2 $T=7820 46240 1 0 $X=7630 $Y=43280
X579 VSS 20 sky130_fd_sc_hd__diode_2 $T=7820 111520 0 0 $X=7630 $Y=111280
X580 VSS 32 sky130_fd_sc_hd__diode_2 $T=7820 155040 0 0 $X=7630 $Y=154800
X581 VSS 34 sky130_fd_sc_hd__diode_2 $T=7820 198560 1 0 $X=7630 $Y=195600
X582 VSS 115 sky130_fd_sc_hd__diode_2 $T=19780 204000 0 0 $X=19590 $Y=203760
X583 VSS 120 sky130_fd_sc_hd__diode_2 $T=23920 111520 0 0 $X=23730 $Y=111280
X584 VSS SCAN_IN<21> sky130_fd_sc_hd__diode_2 $T=34960 176800 0 0 $X=34770 $Y=176560
X585 VSS 215 sky130_fd_sc_hd__diode_2 $T=36340 176800 1 0 $X=36150 $Y=173840
X586 VSS 253 sky130_fd_sc_hd__diode_2 $T=43240 155040 0 0 $X=43050 $Y=154800
X587 VSS 194 sky130_fd_sc_hd__diode_2 $T=47840 100640 0 0 $X=47650 $Y=100400
X588 VSS 337 sky130_fd_sc_hd__diode_2 $T=60260 160480 1 0 $X=60070 $Y=157520
X589 VSS 316 sky130_fd_sc_hd__diode_2 $T=61640 155040 1 0 $X=61450 $Y=152080
X590 VSS 348 sky130_fd_sc_hd__diode_2 $T=68080 182240 0 0 $X=67890 $Y=182000
X591 VSS 378 sky130_fd_sc_hd__diode_2 $T=68540 204000 0 0 $X=68350 $Y=203760
X592 VSS 343 sky130_fd_sc_hd__diode_2 $T=89240 204000 1 0 $X=89050 $Y=201040
X593 VSS 488 sky130_fd_sc_hd__diode_2 $T=92460 127840 1 0 $X=92270 $Y=124880
X594 VSS 507 sky130_fd_sc_hd__diode_2 $T=95220 209440 0 0 $X=95030 $Y=209200
X595 VSS 508 sky130_fd_sc_hd__diode_2 $T=95680 24480 0 0 $X=95490 $Y=24240
X596 VSS SCAN_IN<19> sky130_fd_sc_hd__diode_2 $T=97060 122400 0 0 $X=96870 $Y=122160
X597 VSS 484 sky130_fd_sc_hd__diode_2 $T=98440 187680 0 0 $X=98250 $Y=187440
X598 VSS SCAN_IN<10> sky130_fd_sc_hd__diode_2 $T=99820 57120 0 0 $X=99630 $Y=56880
X599 VSS 585 sky130_fd_sc_hd__diode_2 $T=108560 127840 1 0 $X=108370 $Y=124880
X600 VSS 525 sky130_fd_sc_hd__diode_2 $T=109480 19040 1 0 $X=109290 $Y=16080
X601 VSS 639 sky130_fd_sc_hd__diode_2 $T=120060 89760 1 0 $X=119870 $Y=86800
X602 VSS 568 sky130_fd_sc_hd__diode_2 $T=120060 182240 1 0 $X=119870 $Y=179280
X603 VSS 393 sky130_fd_sc_hd__diode_2 $T=121900 111520 0 0 $X=121710 $Y=111280
X604 VSS 20 sky130_fd_sc_hd__diode_2 $T=121900 144160 0 0 $X=121710 $Y=143920
X605 VSS 20 sky130_fd_sc_hd__diode_2 $T=124660 89760 0 0 $X=124470 $Y=89520
X606 VSS 722 sky130_fd_sc_hd__diode_2 $T=138920 122400 1 0 $X=138730 $Y=119440
X607 VSS 762 sky130_fd_sc_hd__diode_2 $T=145820 19040 1 0 $X=145630 $Y=16080
X608 VSS 674 sky130_fd_sc_hd__diode_2 $T=149040 35360 1 0 $X=148850 $Y=32400
X609 VSS 788 sky130_fd_sc_hd__diode_2 $T=151340 40800 0 0 $X=151150 $Y=40560
X610 VSS 511 sky130_fd_sc_hd__diode_2 $T=154560 89760 0 0 $X=154370 $Y=89520
X611 VSS 530 sky130_fd_sc_hd__diode_2 $T=158700 111520 0 0 $X=158510 $Y=111280
X612 VSS SCAN_IN<0> sky130_fd_sc_hd__diode_2 $T=160540 204000 0 0 $X=160350 $Y=203760
X613 VSS 574 sky130_fd_sc_hd__diode_2 $T=167900 95200 1 0 $X=167710 $Y=92240
X614 VSS 919 sky130_fd_sc_hd__diode_2 $T=178940 89760 0 0 $X=178750 $Y=89520
X615 VSS 712 sky130_fd_sc_hd__diode_2 $T=179400 116960 0 0 $X=179210 $Y=116720
X616 VSS 895 sky130_fd_sc_hd__diode_2 $T=183540 176800 0 0 $X=183350 $Y=176560
X617 VSS 892 sky130_fd_sc_hd__diode_2 $T=184000 127840 0 0 $X=183810 $Y=127600
X618 VSS 950 sky130_fd_sc_hd__diode_2 $T=192280 84320 1 0 $X=192090 $Y=81360
X619 VSS 757 sky130_fd_sc_hd__diode_2 $T=193200 122400 1 0 $X=193010 $Y=119440
X620 VSS 727 sky130_fd_sc_hd__diode_2 $T=194120 149600 1 0 $X=193930 $Y=146640
X621 VSS 961 sky130_fd_sc_hd__diode_2 $T=194580 193120 1 0 $X=194390 $Y=190160
X622 VSS 958 sky130_fd_sc_hd__diode_2 $T=200100 46240 1 0 $X=199910 $Y=43280
X623 VSS 1010 sky130_fd_sc_hd__diode_2 $T=202400 214880 1 0 $X=202210 $Y=211920
X624 VSS 20 sky130_fd_sc_hd__diode_2 $T=205620 122400 0 0 $X=205430 $Y=122160
X625 VSS 1022 sky130_fd_sc_hd__diode_2 $T=206080 116960 1 0 $X=205890 $Y=114000
X626 VSS 996 sky130_fd_sc_hd__diode_2 $T=206540 84320 0 0 $X=206350 $Y=84080
X627 VSS 1007 sky130_fd_sc_hd__diode_2 $T=206540 193120 0 0 $X=206350 $Y=192880
X628 VSS 1040 sky130_fd_sc_hd__diode_2 $T=210220 24480 0 0 $X=210030 $Y=24240
X629 VSS 963 sky130_fd_sc_hd__diode_2 $T=211140 62560 0 0 $X=210950 $Y=62320
X630 VSS VDD 20 ICV_6 $T=7820 209440 1 0 $X=7630 $Y=206480
X631 VSS VDD 54 ICV_6 $T=9660 40800 1 0 $X=9470 $Y=37840
X632 VSS VDD 12 ICV_6 $T=11960 133280 1 0 $X=11770 $Y=130320
X633 VSS VDD 14 ICV_6 $T=12880 144160 1 0 $X=12690 $Y=141200
X634 VSS VDD 73 ICV_6 $T=14260 62560 0 0 $X=14070 $Y=62320
X635 VSS VDD 62 ICV_6 $T=14720 35360 0 0 $X=14530 $Y=35120
X636 VSS VDD 10 ICV_6 $T=21160 95200 1 0 $X=20970 $Y=92240
X637 VSS VDD 171 ICV_6 $T=27600 73440 0 0 $X=27410 $Y=73200
X638 VSS VDD 120 ICV_6 $T=28980 95200 0 0 $X=28790 $Y=94960
X639 VSS VDD 193 ICV_6 $T=34040 57120 1 0 $X=33850 $Y=54160
X640 VSS VDD 92 ICV_6 $T=34040 209440 1 0 $X=33850 $Y=206480
X641 VSS VDD 136 ICV_6 $T=37720 144160 1 0 $X=37530 $Y=141200
X642 VSS VDD 187 ICV_6 $T=38180 155040 1 0 $X=37990 $Y=152080
X643 VSS VDD 228 ICV_6 $T=40020 133280 0 0 $X=39830 $Y=133040
X644 VSS VDD 127 ICV_6 $T=41860 209440 0 0 $X=41670 $Y=209200
X645 VSS VDD 226 ICV_6 $T=42320 100640 0 0 $X=42130 $Y=100400
X646 VSS VDD 279 ICV_6 $T=50140 13600 0 0 $X=49950 $Y=13360
X647 VSS VDD 281 ICV_6 $T=51520 138720 0 0 $X=51330 $Y=138480
X648 VSS VDD 303 ICV_6 $T=54740 35360 1 0 $X=54550 $Y=32400
X649 VSS VDD 17 ICV_6 $T=54740 100640 0 0 $X=54550 $Y=100400
X650 VSS VDD 311 ICV_6 $T=56120 187680 0 0 $X=55930 $Y=187440
X651 VSS VDD 347 ICV_6 $T=62560 144160 1 0 $X=62370 $Y=141200
X652 VSS VDD 312 ICV_6 $T=63020 24480 0 0 $X=62830 $Y=24240
X653 VSS VDD 20 ICV_6 $T=63020 111520 1 0 $X=62830 $Y=108560
X654 VSS VDD 272 ICV_6 $T=65320 209440 0 0 $X=65130 $Y=209200
X655 VSS VDD 351 ICV_6 $T=70380 51680 0 0 $X=70190 $Y=51440
X656 VSS VDD 324 ICV_6 $T=70380 138720 1 0 $X=70190 $Y=135760
X657 VSS VDD 240 ICV_6 $T=70380 204000 1 0 $X=70190 $Y=201040
X658 VSS VDD 393 ICV_6 $T=70840 89760 1 0 $X=70650 $Y=86800
X659 VSS VDD 212 ICV_6 $T=70840 95200 1 0 $X=70650 $Y=92240
X660 VSS VDD 281 ICV_6 $T=71300 95200 0 0 $X=71110 $Y=94960
X661 VSS VDD 378 ICV_6 $T=71300 193120 1 0 $X=71110 $Y=190160
X662 VSS VDD 397 ICV_6 $T=77280 29920 1 0 $X=77090 $Y=26960
X663 VSS VDD 7 ICV_6 $T=79120 106080 1 0 $X=78930 $Y=103120
X664 VSS VDD 400 ICV_6 $T=82340 149600 1 0 $X=82150 $Y=146640
X665 VSS VDD SCAN_IN<7> ICV_6 $T=82800 13600 0 0 $X=82610 $Y=13360
X666 VSS VDD 439 ICV_6 $T=83720 111520 0 0 $X=83530 $Y=111280
X667 VSS VDD 433 ICV_6 $T=84180 176800 1 0 $X=83990 $Y=173840
X668 VSS VDD SCAN_IN<9> ICV_6 $T=91080 24480 0 0 $X=90890 $Y=24240
X669 VSS VDD 473 ICV_6 $T=91080 73440 0 0 $X=90890 $Y=73200
X670 VSS VDD 94 ICV_6 $T=91080 111520 0 0 $X=90890 $Y=111280
X671 VSS VDD 442 ICV_6 $T=91540 225760 1 0 $X=91350 $Y=222800
X672 VSS VDD 144 ICV_6 $T=93380 57120 1 0 $X=93190 $Y=54160
X673 VSS VDD 476 ICV_6 $T=94760 149600 1 0 $X=94570 $Y=146640
X674 VSS VDD 240 ICV_6 $T=97060 209440 1 0 $X=96870 $Y=206480
X675 VSS VDD 520 ICV_6 $T=98900 73440 1 0 $X=98710 $Y=70480
X676 VSS VDD 521 ICV_6 $T=98900 78880 1 0 $X=98710 $Y=75920
X677 VSS VDD 20 ICV_6 $T=99360 29920 1 0 $X=99170 $Y=26960
X678 VSS VDD 523 ICV_6 $T=99360 35360 1 0 $X=99170 $Y=32400
X679 VSS VDD 50 ICV_6 $T=106720 13600 1 0 $X=106530 $Y=10640
X680 VSS VDD 189 ICV_6 $T=109940 182240 0 0 $X=109750 $Y=182000
X681 VSS VDD 582 ICV_6 $T=109940 214880 0 0 $X=109750 $Y=214640
X682 VSS VDD 547 ICV_6 $T=110400 193120 0 0 $X=110210 $Y=192880
X683 VSS VDD 562 ICV_6 $T=115000 89760 1 0 $X=114810 $Y=86800
X684 VSS VDD 190 ICV_6 $T=118220 198560 1 0 $X=118030 $Y=195600
X685 VSS VDD 481 ICV_6 $T=119140 171360 0 0 $X=118950 $Y=171120
X686 VSS VDD 605 ICV_6 $T=121440 127840 1 0 $X=121250 $Y=124880
X687 VSS VDD 641 ICV_6 $T=122820 198560 1 0 $X=122630 $Y=195600
X688 VSS VDD 672 ICV_6 $T=126500 106080 1 0 $X=126310 $Y=103120
X689 VSS VDD 449 ICV_6 $T=126500 111520 1 0 $X=126310 $Y=108560
X690 VSS VDD 555 ICV_6 $T=126500 133280 0 0 $X=126310 $Y=133040
X691 VSS VDD 669 ICV_6 $T=126960 89760 1 0 $X=126770 $Y=86800
X692 VSS VDD 456 ICV_6 $T=126960 95200 1 0 $X=126770 $Y=92240
X693 VSS VDD 659 ICV_6 $T=126960 122400 1 0 $X=126770 $Y=119440
X694 VSS VDD 694 ICV_6 $T=133400 35360 1 0 $X=133210 $Y=32400
X695 VSS VDD 704 ICV_6 $T=133400 100640 1 0 $X=133210 $Y=97680
X696 VSS VDD 700 ICV_6 $T=140760 19040 1 0 $X=140570 $Y=16080
X697 VSS VDD 749 ICV_6 $T=144900 78880 1 0 $X=144710 $Y=75920
X698 VSS VDD 769 ICV_6 $T=147200 144160 0 0 $X=147010 $Y=143920
X699 VSS VDD 767 ICV_6 $T=149500 89760 0 0 $X=149310 $Y=89520
X700 VSS VDD 753 ICV_6 $T=154560 122400 0 0 $X=154370 $Y=122160
X701 VSS VDD 677 ICV_6 $T=155020 73440 0 0 $X=154830 $Y=73200
X702 VSS VDD 563 ICV_6 $T=161460 220320 1 0 $X=161270 $Y=217360
X703 VSS VDD 809 ICV_6 $T=164220 24480 0 0 $X=164030 $Y=24240
X704 VSS VDD 745 ICV_6 $T=167440 138720 0 0 $X=167250 $Y=138480
X705 VSS VDD 883 ICV_6 $T=170200 193120 1 0 $X=170010 $Y=190160
X706 VSS VDD 769 ICV_6 $T=175260 144160 0 0 $X=175070 $Y=143920
X707 VSS VDD 790 ICV_6 $T=175720 116960 1 0 $X=175530 $Y=114000
X708 VSS VDD 906 ICV_6 $T=180320 35360 1 0 $X=180130 $Y=32400
X709 VSS VDD 823 ICV_6 $T=182160 204000 0 0 $X=181970 $Y=203760
X710 VSS VDD 634 ICV_6 $T=182160 220320 1 0 $X=181970 $Y=217360
X711 VSS VDD 20 ICV_6 $T=183540 29920 1 0 $X=183350 $Y=26960
X712 VSS VDD 902 ICV_6 $T=183540 57120 1 0 $X=183350 $Y=54160
X713 VSS VDD 771 ICV_6 $T=183540 95200 1 0 $X=183350 $Y=92240
X714 VSS VDD 952 ICV_6 $T=188600 214880 0 0 $X=188410 $Y=214640
X715 VSS VDD 953 ICV_6 $T=189520 24480 1 0 $X=189330 $Y=21520
X716 VSS VDD 759 ICV_6 $T=189520 138720 0 0 $X=189330 $Y=138480
X717 VSS VDD 947 ICV_6 $T=189520 193120 1 0 $X=189330 $Y=190160
X718 VSS VDD 855 ICV_6 $T=189520 220320 1 0 $X=189330 $Y=217360
X719 VSS VDD 946 ICV_6 $T=190440 187680 0 0 $X=190250 $Y=187440
X720 VSS VDD 948 ICV_6 $T=193660 209440 1 0 $X=193470 $Y=206480
X721 VSS VDD 795 ICV_6 $T=195960 209440 0 0 $X=195770 $Y=209200
X722 VSS VDD 978 ICV_6 $T=203320 160480 0 0 $X=203130 $Y=160240
X723 VSS VDD 1014 ICV_6 $T=210680 209440 1 0 $X=210490 $Y=206480
X724 VSS VDD 1014 ICV_6 $T=210680 214880 1 0 $X=210490 $Y=211920
X725 VSS VDD 1015 ICV_6 $T=211140 111520 1 0 $X=210950 $Y=108560
X726 VSS VDD 1035 ICV_6 $T=216200 116960 0 0 $X=216010 $Y=116720
X727 VSS VDD 1033 ICV_6 $T=216660 198560 0 0 $X=216470 $Y=198320
X728 VSS VDD ICV_7 $T=25760 155040 1 0 $X=25570 $Y=152080
X729 VSS VDD ICV_7 $T=28520 144160 0 0 $X=28330 $Y=143920
X730 VSS VDD ICV_7 $T=28980 214880 1 0 $X=28790 $Y=211920
X731 VSS VDD ICV_7 $T=31280 138720 1 0 $X=31090 $Y=135760
X732 VSS VDD ICV_7 $T=31280 204000 1 0 $X=31090 $Y=201040
X733 VSS VDD ICV_7 $T=41400 182240 0 0 $X=41210 $Y=182000
X734 VSS VDD ICV_7 $T=65780 29920 0 0 $X=65590 $Y=29680
X735 VSS VDD ICV_7 $T=69460 160480 0 0 $X=69270 $Y=160240
X736 VSS VDD ICV_7 $T=76360 204000 0 0 $X=76170 $Y=203760
X737 VSS VDD ICV_7 $T=76360 209440 1 0 $X=76170 $Y=206480
X738 VSS VDD ICV_7 $T=76820 40800 0 0 $X=76630 $Y=40560
X739 VSS VDD ICV_7 $T=84640 84320 0 0 $X=84450 $Y=84080
X740 VSS VDD ICV_7 $T=84640 95200 0 0 $X=84450 $Y=94960
X741 VSS VDD ICV_7 $T=88320 73440 1 0 $X=88130 $Y=70480
X742 VSS VDD ICV_7 $T=95220 187680 1 0 $X=95030 $Y=184720
X743 VSS VDD ICV_7 $T=98900 220320 1 0 $X=98710 $Y=217360
X744 VSS VDD ICV_7 $T=115460 73440 1 0 $X=115270 $Y=70480
X745 VSS VDD ICV_7 $T=123740 13600 0 0 $X=123550 $Y=13360
X746 VSS VDD ICV_7 $T=126960 160480 1 0 $X=126770 $Y=157520
X747 VSS VDD ICV_7 $T=140760 149600 0 0 $X=140570 $Y=149360
X748 VSS VDD ICV_7 $T=166060 57120 1 0 $X=165870 $Y=54160
X749 VSS VDD ICV_7 $T=166060 171360 1 0 $X=165870 $Y=168400
X750 VSS VDD ICV_7 $T=170660 204000 1 0 $X=170470 $Y=201040
X751 VSS VDD ICV_7 $T=183080 68000 1 0 $X=182890 $Y=65040
X752 VSS VDD ICV_7 $T=183080 111520 1 0 $X=182890 $Y=108560
X753 VSS VDD ICV_7 $T=183080 165920 1 0 $X=182890 $Y=162960
X754 VSS VDD ICV_7 $T=198720 78880 1 0 $X=198530 $Y=75920
X755 VSS VDD ICV_7 $T=207920 40800 1 0 $X=207730 $Y=37840
X756 VSS VDD ICV_7 $T=211140 84320 1 0 $X=210950 $Y=81360
X757 VSS VDD ICV_7 $T=211140 171360 1 0 $X=210950 $Y=168400
X758 VSS VDD ICV_7 $T=216660 24480 1 0 $X=216470 $Y=21520
X759 VSS VDD ICV_7 $T=216660 35360 1 0 $X=216470 $Y=32400
X760 VSS VDD ICV_7 $T=216660 35360 0 0 $X=216470 $Y=35120
X761 VSS VDD ICV_7 $T=216660 46240 1 0 $X=216470 $Y=43280
X762 VSS VDD ICV_7 $T=216660 57120 1 0 $X=216470 $Y=54160
X763 VSS VDD ICV_7 $T=216660 89760 1 0 $X=216470 $Y=86800
X764 VSS VDD ICV_7 $T=216660 122400 1 0 $X=216470 $Y=119440
X765 VSS VDD ICV_7 $T=216660 144160 1 0 $X=216470 $Y=141200
X766 VSS VDD ICV_7 $T=216660 149600 1 0 $X=216470 $Y=146640
X767 VSS VDD ICV_7 $T=216660 155040 1 0 $X=216470 $Y=152080
X768 VSS VDD ICV_7 $T=216660 160480 1 0 $X=216470 $Y=157520
X769 VSS VDD ICV_7 $T=216660 165920 1 0 $X=216470 $Y=162960
X770 VSS VDD ICV_7 $T=216660 182240 1 0 $X=216470 $Y=179280
X771 VSS VDD ICV_7 $T=216660 187680 1 0 $X=216470 $Y=184720
X772 VSS VDD ICV_8 $T=117760 127840 0 0 $X=117570 $Y=127600
X773 VSS VDD ICV_8 $T=162380 13600 1 0 $X=162190 $Y=10640
X774 VSS VDD ICV_8 $T=216200 29920 1 0 $X=216010 $Y=26960
X775 VSS VDD ICV_8 $T=216200 40800 1 0 $X=216010 $Y=37840
X776 VSS VDD ICV_8 $T=216200 62560 1 0 $X=216010 $Y=59600
X777 VSS VDD ICV_8 $T=216200 68000 1 0 $X=216010 $Y=65040
X778 VSS VDD ICV_8 $T=216200 84320 1 0 $X=216010 $Y=81360
X779 VSS VDD ICV_8 $T=216200 95200 1 0 $X=216010 $Y=92240
X780 VSS VDD ICV_8 $T=216200 106080 1 0 $X=216010 $Y=103120
X781 VSS VDD ICV_8 $T=216200 111520 1 0 $X=216010 $Y=108560
X782 VSS VDD ICV_8 $T=216200 116960 1 0 $X=216010 $Y=114000
X783 VSS VDD ICV_8 $T=216200 127840 1 0 $X=216010 $Y=124880
X784 VSS VDD ICV_8 $T=216200 133280 1 0 $X=216010 $Y=130320
X785 VSS VDD ICV_8 $T=216200 171360 1 0 $X=216010 $Y=168400
X786 VSS VDD ICV_8 $T=216200 198560 1 0 $X=216010 $Y=195600
X787 VSS VDD ICV_8 $T=216200 209440 1 0 $X=216010 $Y=206480
X788 VSS VDD ICV_8 $T=216200 214880 1 0 $X=216010 $Y=211920
X789 VSS VDD ICV_8 $T=216200 220320 1 0 $X=216010 $Y=217360
X790 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 35360 0 0 $X=6710 $Y=35120
X791 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 209440 0 0 $X=6710 $Y=209200
X792 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=14260 149600 1 0 $X=14070 $Y=146640
X793 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=14260 155040 1 0 $X=14070 $Y=152080
X794 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=20240 111520 1 0 $X=20050 $Y=108560
X795 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=25300 89760 1 0 $X=25110 $Y=86800
X796 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=33120 111520 1 0 $X=32930 $Y=108560
X797 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=38180 95200 1 0 $X=37990 $Y=92240
X798 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=40480 24480 1 0 $X=40290 $Y=21520
X799 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=40480 40800 1 0 $X=40290 $Y=37840
X800 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=40480 182240 1 0 $X=40290 $Y=179280
X801 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=42320 176800 1 0 $X=42130 $Y=173840
X802 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=53360 51680 1 0 $X=53170 $Y=48720
X803 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=54280 95200 1 0 $X=54090 $Y=92240
X804 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=54740 182240 1 0 $X=54550 $Y=179280
X805 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=56580 225760 1 0 $X=56390 $Y=222800
X806 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=59800 138720 1 0 $X=59610 $Y=135760
X807 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=61640 214880 1 0 $X=61450 $Y=211920
X808 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=62100 106080 1 0 $X=61910 $Y=103120
X809 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=62100 204000 0 0 $X=61910 $Y=203760
X810 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=64400 204000 1 0 $X=64210 $Y=201040
X811 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=68540 149600 1 0 $X=68350 $Y=146640
X812 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69000 40800 1 0 $X=68810 $Y=37840
X813 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69920 160480 1 0 $X=69730 $Y=157520
X814 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=76360 35360 1 0 $X=76170 $Y=32400
X815 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=80960 165920 0 0 $X=80770 $Y=165680
X816 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=84180 155040 1 0 $X=83990 $Y=152080
X817 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=96140 193120 1 0 $X=95950 $Y=190160
X818 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=97980 225760 1 0 $X=97790 $Y=222800
X819 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=102580 138720 0 0 $X=102390 $Y=138480
X820 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=111780 127840 0 0 $X=111590 $Y=127600
X821 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=114540 182240 1 0 $X=114350 $Y=179280
X822 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=115920 95200 1 0 $X=115730 $Y=92240
X823 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=115920 100640 1 0 $X=115730 $Y=97680
X824 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=121900 57120 1 0 $X=121710 $Y=54160
X825 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=122360 138720 0 0 $X=122170 $Y=138480
X826 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=124660 24480 1 0 $X=124470 $Y=21520
X827 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=125580 155040 1 0 $X=125390 $Y=152080
X828 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=125580 204000 1 0 $X=125390 $Y=201040
X829 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=126500 133280 1 0 $X=126310 $Y=130320
X830 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=126500 149600 1 0 $X=126310 $Y=146640
X831 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=126500 209440 1 0 $X=126310 $Y=206480
X832 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=137080 89760 0 0 $X=136890 $Y=89520
X833 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=138920 13600 1 0 $X=138730 $Y=10640
X834 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=138920 51680 1 0 $X=138730 $Y=48720
X835 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=140300 198560 1 0 $X=140110 $Y=195600
X836 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=140760 204000 1 0 $X=140570 $Y=201040
X837 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=141220 106080 1 0 $X=141030 $Y=103120
X838 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146280 155040 1 0 $X=146090 $Y=152080
X839 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146740 225760 1 0 $X=146550 $Y=222800
X840 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=150880 171360 1 0 $X=150690 $Y=168400
X841 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=152720 57120 1 0 $X=152530 $Y=54160
X842 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=152720 62560 1 0 $X=152530 $Y=59600
X843 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=152720 73440 1 0 $X=152530 $Y=70480
X844 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=153640 35360 0 0 $X=153450 $Y=35120
X845 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=153640 111520 1 0 $X=153450 $Y=108560
X846 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=153640 127840 0 0 $X=153450 $Y=127600
X847 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=156400 51680 0 0 $X=156210 $Y=51440
X848 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=160540 155040 0 0 $X=160350 $Y=154800
X849 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=164680 193120 1 0 $X=164490 $Y=190160
X850 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=167440 46240 1 0 $X=167250 $Y=43280
X851 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=167440 106080 0 0 $X=167250 $Y=105840
X852 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=172040 62560 1 0 $X=171850 $Y=59600
X853 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=175260 95200 1 0 $X=175070 $Y=92240
X854 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=177560 68000 1 0 $X=177370 $Y=65040
X855 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=178020 214880 1 0 $X=177830 $Y=211920
X856 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=178940 133280 1 0 $X=178750 $Y=130320
X857 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=181700 84320 1 0 $X=181510 $Y=81360
X858 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=182620 62560 1 0 $X=182430 $Y=59600
X859 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=185380 106080 0 0 $X=185190 $Y=105840
X860 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=187220 155040 0 0 $X=187030 $Y=154800
X861 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=189520 198560 0 0 $X=189330 $Y=198320
X862 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=190900 29920 1 0 $X=190710 $Y=26960
X863 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=197340 171360 1 0 $X=197150 $Y=168400
X864 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=200560 19040 1 0 $X=200370 $Y=16080
X865 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=212980 13600 1 0 $X=212790 $Y=10640
X866 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=215740 13600 0 0 $X=215550 $Y=13360
X867 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=216200 127840 0 0 $X=216010 $Y=127600
X868 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=216200 144160 0 0 $X=216010 $Y=143920
X869 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=216200 176800 0 0 $X=216010 $Y=176560
X870 VSS VDD 16 ICV_9 $T=11040 225760 1 0 $X=10850 $Y=222800
X871 VSS VDD 32 ICV_9 $T=11960 171360 1 0 $X=11770 $Y=168400
X872 VSS VDD 81 ICV_9 $T=13340 57120 1 0 $X=13150 $Y=54160
X873 VSS VDD 116 ICV_9 $T=20700 13600 0 0 $X=20510 $Y=13360
X874 VSS VDD 25 ICV_9 $T=21160 51680 1 0 $X=20970 $Y=48720
X875 VSS VDD 136 ICV_9 $T=34960 122400 0 0 $X=34770 $Y=122160
X876 VSS VDD 233 ICV_9 $T=39560 122400 1 0 $X=39370 $Y=119440
X877 VSS VDD 225 ICV_9 $T=40940 214880 1 0 $X=40750 $Y=211920
X878 VSS VDD 212 ICV_9 $T=41400 19040 1 0 $X=41210 $Y=16080
X879 VSS VDD 240 ICV_9 $T=41400 209440 1 0 $X=41210 $Y=206480
X880 VSS VDD 230 ICV_9 $T=41860 144160 0 0 $X=41670 $Y=143920
X881 VSS VDD 248 ICV_9 $T=48300 144160 0 0 $X=48110 $Y=143920
X882 VSS VDD 231 ICV_9 $T=49220 171360 1 0 $X=49030 $Y=168400
X883 VSS VDD 258 ICV_9 $T=51520 149600 1 0 $X=51330 $Y=146640
X884 VSS VDD 286 ICV_9 $T=54280 182240 0 0 $X=54090 $Y=182000
X885 VSS VDD 307 ICV_9 $T=55200 40800 0 0 $X=55010 $Y=40560
X886 VSS VDD 266 ICV_9 $T=55200 89760 0 0 $X=55010 $Y=89520
X887 VSS VDD 258 ICV_9 $T=63020 160480 0 0 $X=62830 $Y=160240
X888 VSS VDD CLK_OUT ICV_9 $T=63940 89760 1 0 $X=63750 $Y=86800
X889 VSS VDD 364 ICV_9 $T=65780 171360 1 0 $X=65590 $Y=168400
X890 VSS VDD 372 ICV_9 $T=67620 35360 1 0 $X=67430 $Y=32400
X891 VSS VDD 355 ICV_9 $T=68080 127840 0 0 $X=67890 $Y=127600
X892 VSS VDD 359 ICV_9 $T=68540 225760 1 0 $X=68350 $Y=222800
X893 VSS VDD 289 ICV_9 $T=69000 57120 1 0 $X=68810 $Y=54160
X894 VSS VDD 276 ICV_9 $T=77280 73440 0 0 $X=77090 $Y=73200
X895 VSS VDD 417 ICV_9 $T=77280 78880 1 0 $X=77090 $Y=75920
X896 VSS VDD 421 ICV_9 $T=77280 89760 1 0 $X=77090 $Y=86800
X897 VSS VDD 420 ICV_9 $T=80500 220320 0 0 $X=80310 $Y=220080
X898 VSS VDD 416 ICV_9 $T=80960 68000 0 0 $X=80770 $Y=67760
X899 VSS VDD 428 ICV_9 $T=82340 138720 1 0 $X=82150 $Y=135760
X900 VSS VDD 459 ICV_9 $T=91080 187680 0 0 $X=90890 $Y=187440
X901 VSS VDD 17 ICV_9 $T=93380 68000 0 0 $X=93190 $Y=67760
X902 VSS VDD 20 ICV_9 $T=93840 62560 1 0 $X=93650 $Y=59600
X903 VSS VDD 496 ICV_9 $T=93840 68000 1 0 $X=93650 $Y=65040
X904 VSS VDD 377 ICV_9 $T=93840 149600 0 0 $X=93650 $Y=149360
X905 VSS VDD 473 ICV_9 $T=95680 100640 1 0 $X=95490 $Y=97680
X906 VSS VDD 451 ICV_9 $T=96140 84320 1 0 $X=95950 $Y=81360
X907 VSS VDD 511 ICV_9 $T=96600 95200 1 0 $X=96410 $Y=92240
X908 VSS VDD 245 ICV_9 $T=97060 214880 1 0 $X=96870 $Y=211920
X909 VSS VDD 473 ICV_9 $T=98440 78880 0 0 $X=98250 $Y=78640
X910 VSS VDD 521 ICV_9 $T=105340 46240 1 0 $X=105150 $Y=43280
X911 VSS VDD 130 ICV_9 $T=105340 57120 1 0 $X=105150 $Y=54160
X912 VSS VDD 586 ICV_9 $T=111320 13600 1 0 $X=111130 $Y=10640
X913 VSS VDD 566 ICV_9 $T=111320 84320 1 0 $X=111130 $Y=81360
X914 VSS VDD 597 ICV_9 $T=111320 95200 0 0 $X=111130 $Y=94960
X915 VSS VDD 599 ICV_9 $T=111320 106080 0 0 $X=111130 $Y=105840
X916 VSS VDD 537 ICV_9 $T=111780 133280 1 0 $X=111590 $Y=130320
X917 VSS VDD 301 ICV_9 $T=117760 214880 1 0 $X=117570 $Y=211920
X918 VSS VDD 529 ICV_9 $T=120060 62560 1 0 $X=119870 $Y=59600
X919 VSS VDD 630 ICV_9 $T=121440 138720 1 0 $X=121250 $Y=135760
X920 VSS VDD 548 ICV_9 $T=123740 116960 1 0 $X=123550 $Y=114000
X921 VSS VDD 667 ICV_9 $T=124660 165920 1 0 $X=124470 $Y=162960
X922 VSS VDD 656 ICV_9 $T=128340 95200 0 0 $X=128150 $Y=94960
X923 VSS VDD 666 ICV_9 $T=132480 51680 0 0 $X=132290 $Y=51440
X924 VSS VDD 718 ICV_9 $T=136160 149600 1 0 $X=135970 $Y=146640
X925 VSS VDD 678 ICV_9 $T=137540 155040 0 0 $X=137350 $Y=154800
X926 VSS VDD 725 ICV_9 $T=139380 24480 0 0 $X=139190 $Y=24240
X927 VSS VDD 509 ICV_9 $T=143060 144160 1 0 $X=142870 $Y=141200
X928 VSS VDD 744 ICV_9 $T=149500 46240 0 0 $X=149310 $Y=46000
X929 VSS VDD 752 ICV_9 $T=149500 171360 0 0 $X=149310 $Y=171120
X930 VSS VDD 726 ICV_9 $T=149960 100640 1 0 $X=149770 $Y=97680
X931 VSS VDD 766 ICV_9 $T=151340 68000 1 0 $X=151150 $Y=65040
X932 VSS VDD 325 ICV_9 $T=151800 165920 1 0 $X=151610 $Y=162960
X933 VSS VDD 325 ICV_9 $T=155940 160480 0 0 $X=155750 $Y=160240
X934 VSS VDD 798 ICV_9 $T=159160 193120 0 0 $X=158970 $Y=192880
X935 VSS VDD 864 ICV_9 $T=167900 13600 1 0 $X=167710 $Y=10640
X936 VSS VDD 901 ICV_9 $T=175260 209440 0 0 $X=175070 $Y=209200
X937 VSS VDD 765 ICV_9 $T=176180 62560 0 0 $X=175990 $Y=62320
X938 VSS VDD 853 ICV_9 $T=178020 13600 1 0 $X=177830 $Y=10640
X939 VSS VDD 927 ICV_9 $T=180780 89760 1 0 $X=180590 $Y=86800
X940 VSS VDD 930 ICV_9 $T=181700 40800 1 0 $X=181510 $Y=37840
X941 VSS VDD 830 ICV_9 $T=187220 19040 0 0 $X=187030 $Y=18800
X942 VSS VDD 932 ICV_9 $T=192280 95200 1 0 $X=192090 $Y=92240
X943 VSS VDD 967 ICV_9 $T=193660 122400 0 0 $X=193470 $Y=122160
X944 VSS VDD 987 ICV_9 $T=201020 106080 1 0 $X=200830 $Y=103120
X945 VSS VDD 928 ICV_9 $T=203320 144160 0 0 $X=203130 $Y=143920
X946 VSS VDD 844 ICV_9 $T=207460 106080 0 0 $X=207270 $Y=105840
X947 VSS VDD 995 ICV_9 $T=208380 89760 1 0 $X=208190 $Y=86800
X948 VSS VDD 1039 ICV_9 $T=213900 133280 0 0 $X=213710 $Y=133040
X949 VSS VDD 1044 ICV_9 $T=214360 171360 0 0 $X=214170 $Y=171120
X950 VSS VDD 1038 ICV_9 $T=215280 73440 0 0 $X=215090 $Y=73200
X951 VSS VDD ICV_10 $T=18400 127840 1 0 $X=18210 $Y=124880
X952 VSS VDD ICV_10 $T=18400 171360 1 0 $X=18210 $Y=168400
X953 VSS VDD ICV_10 $T=18400 220320 1 0 $X=18210 $Y=217360
X954 VSS VDD ICV_10 $T=32200 73440 0 0 $X=32010 $Y=73200
X955 VSS VDD ICV_10 $T=32200 116960 0 0 $X=32010 $Y=116720
X956 VSS VDD ICV_10 $T=46460 73440 1 0 $X=46270 $Y=70480
X957 VSS VDD ICV_10 $T=46920 13600 1 0 $X=46730 $Y=10640
X958 VSS VDD ICV_10 $T=60260 46240 0 0 $X=60070 $Y=46000
X959 VSS VDD ICV_10 $T=60260 84320 0 0 $X=60070 $Y=84080
X960 VSS VDD ICV_10 $T=60260 160480 0 0 $X=60070 $Y=160240
X961 VSS VDD ICV_10 $T=60260 204000 0 0 $X=60070 $Y=203760
X962 VSS VDD ICV_10 $T=60260 214880 0 0 $X=60070 $Y=214640
X963 VSS VDD ICV_10 $T=74520 40800 1 0 $X=74330 $Y=37840
X964 VSS VDD ICV_10 $T=74520 127840 1 0 $X=74330 $Y=124880
X965 VSS VDD ICV_10 $T=88320 111520 0 0 $X=88130 $Y=111280
X966 VSS VDD ICV_10 $T=102580 19040 1 0 $X=102390 $Y=16080
X967 VSS VDD ICV_10 $T=102580 62560 1 0 $X=102390 $Y=59600
X968 VSS VDD ICV_10 $T=102580 84320 1 0 $X=102390 $Y=81360
X969 VSS VDD ICV_10 $T=102580 138720 1 0 $X=102390 $Y=135760
X970 VSS VDD ICV_10 $T=116380 46240 0 0 $X=116190 $Y=46000
X971 VSS VDD ICV_10 $T=116380 111520 0 0 $X=116190 $Y=111280
X972 VSS VDD ICV_10 $T=116380 171360 0 0 $X=116190 $Y=171120
X973 VSS VDD ICV_10 $T=144440 133280 0 0 $X=144250 $Y=133040
X974 VSS VDD ICV_10 $T=144440 204000 0 0 $X=144250 $Y=203760
X975 VSS VDD ICV_10 $T=144440 209440 0 0 $X=144250 $Y=209200
X976 VSS VDD ICV_10 $T=158700 29920 1 0 $X=158510 $Y=26960
X977 VSS VDD ICV_10 $T=158700 116960 1 0 $X=158510 $Y=114000
X978 VSS VDD ICV_10 $T=172500 40800 0 0 $X=172310 $Y=40560
X979 VSS VDD ICV_10 $T=186760 127840 1 0 $X=186570 $Y=124880
X980 VSS VDD ICV_10 $T=186760 133280 1 0 $X=186570 $Y=130320
X981 VSS VDD ICV_10 $T=186760 155040 1 0 $X=186570 $Y=152080
X982 VSS VDD ICV_10 $T=186760 220320 1 0 $X=186570 $Y=217360
X983 VSS VDD ICV_10 $T=200560 138720 0 0 $X=200370 $Y=138480
X984 VSS VDD ICV_10 $T=200560 160480 0 0 $X=200370 $Y=160240
X985 VSS VDD ICV_10 $T=200560 209440 0 0 $X=200370 $Y=209200
X986 VSS VDD ICV_10 $T=214820 57120 1 0 $X=214630 $Y=54160
X987 VSS VDD ICV_10 $T=214820 89760 1 0 $X=214630 $Y=86800
X988 VSS VDD ICV_10 $T=214820 144160 1 0 $X=214630 $Y=141200
X989 VSS VDD ICV_10 $T=214820 149600 1 0 $X=214630 $Y=146640
X990 VSS VDD ICV_10 $T=214820 165920 1 0 $X=214630 $Y=162960
X991 VSS VDD ICV_11 $T=11960 13600 1 0 $X=11770 $Y=10640
X992 VSS VDD ICV_11 $T=12420 209440 0 0 $X=12230 $Y=209200
X993 VSS VDD ICV_11 $T=20240 160480 1 0 $X=20050 $Y=157520
X994 VSS VDD ICV_11 $T=25760 84320 0 0 $X=25570 $Y=84080
X995 VSS VDD ICV_11 $T=27600 171360 1 0 $X=27410 $Y=168400
X996 VSS VDD ICV_11 $T=37720 149600 0 0 $X=37530 $Y=149360
X997 VSS VDD ICV_11 $T=53820 165920 0 0 $X=53630 $Y=165680
X998 VSS VDD ICV_11 $T=55660 171360 1 0 $X=55470 $Y=168400
X999 VSS VDD ICV_11 $T=62100 13600 0 0 $X=61910 $Y=13360
X1000 VSS VDD ICV_11 $T=75900 193120 0 0 $X=75710 $Y=192880
X1001 VSS VDD ICV_11 $T=90160 19040 0 0 $X=89970 $Y=18800
X1002 VSS VDD ICV_11 $T=103500 106080 0 0 $X=103310 $Y=105840
X1003 VSS VDD ICV_11 $T=111780 138720 1 0 $X=111590 $Y=135760
X1004 VSS VDD ICV_11 $T=124200 214880 1 0 $X=124010 $Y=211920
X1005 VSS VDD ICV_11 $T=128800 165920 0 0 $X=128610 $Y=165680
X1006 VSS VDD ICV_11 $T=132480 62560 1 0 $X=132290 $Y=59600
X1007 VSS VDD ICV_11 $T=138000 176800 1 0 $X=137810 $Y=173840
X1008 VSS VDD ICV_11 $T=138460 68000 0 0 $X=138270 $Y=67760
X1009 VSS VDD ICV_11 $T=147200 116960 1 0 $X=147010 $Y=114000
X1010 VSS VDD ICV_11 $T=152260 225760 1 0 $X=152070 $Y=222800
X1011 VSS VDD ICV_11 $T=166520 138720 1 0 $X=166330 $Y=135760
X1012 VSS VDD ICV_11 $T=172500 171360 1 0 $X=172310 $Y=168400
X1013 VSS VDD ICV_11 $T=180320 198560 1 0 $X=180130 $Y=195600
X1014 VSS VDD ICV_11 $T=182160 78880 0 0 $X=181970 $Y=78640
X1015 VSS VDD ICV_11 $T=208380 68000 1 0 $X=208190 $Y=65040
X1016 VSS VDD ICV_11 $T=213900 46240 0 0 $X=213710 $Y=46000
X1017 VSS VDD ICV_11 $T=213900 106080 0 0 $X=213710 $Y=105840
X1018 VSS VDD ICV_11 $T=214360 78880 0 0 $X=214170 $Y=78640
X1019 VSS VDD ICV_11 $T=214360 138720 0 0 $X=214170 $Y=138480
X1020 VSS VDD ICV_11 $T=214360 214880 0 0 $X=214170 $Y=214640
X1021 VSS VDD ICV_12 $T=17940 24480 1 0 $X=17750 $Y=21520
X1022 VSS VDD ICV_12 $T=17940 111520 1 0 $X=17750 $Y=108560
X1023 VSS VDD ICV_12 $T=17940 116960 1 0 $X=17750 $Y=114000
X1024 VSS VDD ICV_12 $T=17940 122400 1 0 $X=17750 $Y=119440
X1025 VSS VDD ICV_12 $T=17940 214880 1 0 $X=17750 $Y=211920
X1026 VSS VDD ICV_12 $T=17940 225760 0 0 $X=17750 $Y=225520
X1027 VSS VDD ICV_12 $T=31740 51680 0 0 $X=31550 $Y=51440
X1028 VSS VDD ICV_12 $T=46000 24480 1 0 $X=45810 $Y=21520
X1029 VSS VDD ICV_12 $T=46000 29920 1 0 $X=45810 $Y=26960
X1030 VSS VDD ICV_12 $T=46000 40800 1 0 $X=45810 $Y=37840
X1031 VSS VDD ICV_12 $T=46000 116960 1 0 $X=45810 $Y=114000
X1032 VSS VDD ICV_12 $T=46000 122400 1 0 $X=45810 $Y=119440
X1033 VSS VDD ICV_12 $T=46000 155040 1 0 $X=45810 $Y=152080
X1034 VSS VDD ICV_12 $T=46000 182240 1 0 $X=45810 $Y=179280
X1035 VSS VDD ICV_12 $T=59800 106080 0 0 $X=59610 $Y=105840
X1036 VSS VDD ICV_12 $T=74060 35360 1 0 $X=73870 $Y=32400
X1037 VSS VDD ICV_12 $T=74060 149600 1 0 $X=73870 $Y=146640
X1038 VSS VDD ICV_12 $T=74060 187680 1 0 $X=73870 $Y=184720
X1039 VSS VDD ICV_12 $T=102120 100640 1 0 $X=101930 $Y=97680
X1040 VSS VDD ICV_12 $T=102120 127840 1 0 $X=101930 $Y=124880
X1041 VSS VDD ICV_12 $T=117760 13600 1 0 $X=117570 $Y=10640
X1042 VSS VDD ICV_12 $T=130180 19040 1 0 $X=129990 $Y=16080
X1043 VSS VDD ICV_12 $T=130180 24480 1 0 $X=129990 $Y=21520
X1044 VSS VDD ICV_12 $T=130180 116960 1 0 $X=129990 $Y=114000
X1045 VSS VDD ICV_12 $T=143980 46240 0 0 $X=143790 $Y=46000
X1046 VSS VDD ICV_12 $T=143980 155040 0 0 $X=143790 $Y=154800
X1047 VSS VDD ICV_12 $T=158240 62560 1 0 $X=158050 $Y=59600
X1048 VSS VDD ICV_12 $T=158240 73440 1 0 $X=158050 $Y=70480
X1049 VSS VDD ICV_12 $T=158240 127840 1 0 $X=158050 $Y=124880
X1050 VSS VDD ICV_12 $T=158240 198560 1 0 $X=158050 $Y=195600
X1051 VSS VDD ICV_12 $T=200100 19040 0 0 $X=199910 $Y=18800
X1052 VSS VDD ICV_12 $T=200100 111520 0 0 $X=199910 $Y=111280
X1053 VSS VDD ICV_12 $T=214360 35360 1 0 $X=214170 $Y=32400
X1054 VSS VDD ICV_12 $T=214360 160480 1 0 $X=214170 $Y=157520
X1055 VSS VDD 59 65 VDD 34 VSS sky130_fd_sc_hd__nor2_4 $T=9660 198560 1 0 $X=9470 $Y=195600
X1056 VSS VDD 61 35 VDD 53 VSS sky130_fd_sc_hd__nor2_4 $T=10120 24480 1 0 $X=9930 $Y=21520
X1057 VSS VDD 25 107 VDD 88 VSS sky130_fd_sc_hd__nor2_4 $T=21160 57120 1 0 $X=20970 $Y=54160
X1058 VSS VDD 118 131 VDD 122 VSS sky130_fd_sc_hd__nor2_4 $T=23460 171360 1 0 $X=23270 $Y=168400
X1059 VSS VDD 61 134 VDD 167 VSS sky130_fd_sc_hd__nor2_4 $T=23920 35360 0 0 $X=23730 $Y=35120
X1060 VSS VDD 120 159 VDD 180 VSS sky130_fd_sc_hd__nor2_4 $T=25760 111520 0 0 $X=25570 $Y=111280
X1061 VSS VDD 172 211 VDD 201 VSS sky130_fd_sc_hd__nor2_4 $T=34040 95200 1 0 $X=33850 $Y=92240
X1062 VSS VDD 191 124 VDD 203 VSS sky130_fd_sc_hd__nor2_4 $T=36340 24480 1 0 $X=36150 $Y=21520
X1063 VSS VDD 173 222 VDD 215 VSS sky130_fd_sc_hd__nor2_4 $T=38180 176800 1 0 $X=37990 $Y=173840
X1064 VSS VDD 128 350 VDD 239 VSS sky130_fd_sc_hd__nor2_4 $T=60720 46240 1 0 $X=60530 $Y=43280
X1065 VSS VDD 307 351 VDD 333 VSS sky130_fd_sc_hd__nor2_4 $T=61640 57120 1 0 $X=61450 $Y=54160
X1066 VSS VDD 147 376 VDD 298 VSS sky130_fd_sc_hd__nor2_4 $T=68080 24480 1 0 $X=67890 $Y=21520
X1067 VSS VDD 370 CLK_OUT VDD 380 VSS sky130_fd_sc_hd__nor2_4 $T=71300 100640 0 0 $X=71110 $Y=100400
X1068 VSS VDD SCAN_IN<18> 315 VDD 438 VSS sky130_fd_sc_hd__nor2_4 $T=77280 111520 0 0 $X=77090 $Y=111280
X1069 VSS VDD 484 145 VDD 546 VSS sky130_fd_sc_hd__nor2_4 $T=100280 187680 0 0 $X=100090 $Y=187440
X1070 VSS VDD 565 562 VDD 536 VSS sky130_fd_sc_hd__nor2_4 $T=109940 89760 0 0 $X=109750 $Y=89520
X1071 VSS VDD 529 591 VDD 572 VSS sky130_fd_sc_hd__nor2_4 $T=115000 62560 1 0 $X=114810 $Y=59600
X1072 VSS VDD 507 549 VDD 610 VSS sky130_fd_sc_hd__nor2_4 $T=115920 165920 1 0 $X=115730 $Y=162960
X1073 VSS VDD 623 655 VDD 603 VSS sky130_fd_sc_hd__nor2_4 $T=120520 24480 1 0 $X=120330 $Y=21520
X1074 VSS VDD 620 625 VDD 617 VSS sky130_fd_sc_hd__nor2_4 $T=122820 160480 1 0 $X=122630 $Y=157520
X1075 VSS VDD SCAN_IN<11> 661 VDD 705 VSS sky130_fd_sc_hd__nor2_4 $T=130180 127840 0 0 $X=129990 $Y=127600
X1076 VSS VDD 696 300 VDD 681 VSS sky130_fd_sc_hd__nor2_4 $T=132020 198560 0 0 $X=131830 $Y=198320
X1077 VSS VDD 511 608 VDD 806 VSS sky130_fd_sc_hd__nor2_4 $T=156400 89760 0 0 $X=156210 $Y=89520
X1078 VSS VDD 889 907 VDD 857 VSS sky130_fd_sc_hd__nor2_4 $T=175720 204000 1 0 $X=175530 $Y=201040
X1079 VSS VDD 924 931 VDD 741 VSS sky130_fd_sc_hd__nor2_4 $T=180320 171360 1 0 $X=180130 $Y=168400
X1080 VSS VDD 952 938 VDD 896 VSS sky130_fd_sc_hd__nor2_4 $T=189520 214880 1 0 $X=189330 $Y=211920
X1081 VSS VDD 1009 970 VDD 974 VSS sky130_fd_sc_hd__nor2_4 $T=203320 78880 0 0 $X=203130 $Y=78640
X1082 VSS VDD 1013 979 VDD 995 VSS sky130_fd_sc_hd__nor2_4 $T=204240 187680 0 0 $X=204050 $Y=187440
X1083 VSS VDD 1024 1036 VDD 1020 VSS sky130_fd_sc_hd__nor2_4 $T=208380 19040 1 0 $X=208190 $Y=16080
X1084 VSS VDD 911 1037 VDD 1045 VSS sky130_fd_sc_hd__nor2_4 $T=212980 40800 0 0 $X=212790 $Y=40560
X1085 VSS VDD 963 1038 VDD 1046 VSS sky130_fd_sc_hd__nor2_4 $T=212980 62560 0 0 $X=212790 $Y=62320
X1086 VSS VDD 1048 1025 VDD 1052 VSS sky130_fd_sc_hd__nor2_4 $T=213900 165920 0 0 $X=213710 $Y=165680
X1087 VSS VDD 24 VDD 11 VSS sky130_fd_sc_hd__inv_8 $T=7820 73440 0 0 $X=7630 $Y=73200
X1088 VSS VDD BB_IN VDD 46 VSS sky130_fd_sc_hd__inv_8 $T=7820 144160 1 0 $X=7630 $Y=141200
X1089 VSS VDD 33 VDD 32 VSS sky130_fd_sc_hd__inv_8 $T=7820 171360 0 0 $X=7630 $Y=171120
X1090 VSS VDD 81 VDD 73 VSS sky130_fd_sc_hd__inv_8 $T=13340 57120 0 0 $X=13150 $Y=56880
X1091 VSS VDD 98 VDD 120 VSS sky130_fd_sc_hd__inv_8 $T=21160 116960 1 0 $X=20970 $Y=114000
X1092 VSS VDD 105 VDD 148 VSS sky130_fd_sc_hd__inv_8 $T=21160 155040 0 0 $X=20970 $Y=154800
X1093 VSS VDD 115 VDD 79 VSS sky130_fd_sc_hd__inv_8 $T=21160 214880 1 0 $X=20970 $Y=211920
X1094 VSS VDD 129 VDD 164 VSS sky130_fd_sc_hd__inv_8 $T=23460 73440 1 0 $X=23270 $Y=70480
X1095 VSS VDD 172 VDD 37 VSS sky130_fd_sc_hd__inv_8 $T=26220 95200 1 0 $X=26030 $Y=92240
X1096 VSS VDD 187 VDD 136 VSS sky130_fd_sc_hd__inv_8 $T=32660 144160 1 0 $X=32470 $Y=141200
X1097 VSS VDD 149 VDD 132 VSS sky130_fd_sc_hd__inv_8 $T=37260 182240 0 0 $X=37070 $Y=182000
X1098 VSS VDD 199 VDD 235 VSS sky130_fd_sc_hd__inv_8 $T=39100 84320 1 0 $X=38910 $Y=81360
X1099 VSS VDD 210 VDD 246 VSS sky130_fd_sc_hd__inv_8 $T=40020 62560 1 0 $X=39830 $Y=59600
X1100 VSS VDD 214 VDD 226 VSS sky130_fd_sc_hd__inv_8 $T=43240 106080 0 0 $X=43050 $Y=105840
X1101 VSS VDD 232 VDD 264 VSS sky130_fd_sc_hd__inv_8 $T=43700 35360 0 0 $X=43510 $Y=35120
X1102 VSS VDD 249 VDD 258 VSS sky130_fd_sc_hd__inv_8 $T=46460 187680 0 0 $X=46270 $Y=187440
X1103 VSS VDD 272 VDD 150 VSS sky130_fd_sc_hd__inv_8 $T=48760 198560 0 0 $X=48570 $Y=198320
X1104 VSS VDD 243 VDD 241 VSS sky130_fd_sc_hd__inv_8 $T=49680 73440 1 0 $X=49490 $Y=70480
X1105 VSS VDD 273 VDD 265 VSS sky130_fd_sc_hd__inv_8 $T=51060 51680 0 0 $X=50870 $Y=51440
X1106 VSS VDD 324 VDD 327 VSS sky130_fd_sc_hd__inv_8 $T=57500 144160 1 0 $X=57310 $Y=141200
X1107 VSS VDD 317 VDD 274 VSS sky130_fd_sc_hd__inv_8 $T=63020 19040 0 0 $X=62830 $Y=18800
X1108 VSS VDD 334 VDD 370 VSS sky130_fd_sc_hd__inv_8 $T=63020 100640 0 0 $X=62830 $Y=100400
X1109 VSS VDD 251 VDD 372 VSS sky130_fd_sc_hd__inv_8 $T=65320 35360 0 0 $X=65130 $Y=35120
X1110 VSS VDD 355 VDD 247 VSS sky130_fd_sc_hd__inv_8 $T=68080 122400 1 0 $X=67890 $Y=119440
X1111 VSS VDD 356 VDD 347 VSS sky130_fd_sc_hd__inv_8 $T=68080 144160 1 0 $X=67890 $Y=141200
X1112 VSS VDD 353 VDD 338 VSS sky130_fd_sc_hd__inv_8 $T=72220 176800 0 0 $X=72030 $Y=176560
X1113 VSS VDD 331 VDD 400 VSS sky130_fd_sc_hd__inv_8 $T=77280 149600 1 0 $X=77090 $Y=146640
X1114 VSS VDD 439 VDD 432 VSS sky130_fd_sc_hd__inv_8 $T=83720 116960 1 0 $X=83530 $Y=114000
X1115 VSS VDD SCAN_IN<19> VDD 413 VSS sky130_fd_sc_hd__inv_8 $T=87860 111520 1 0 $X=87670 $Y=108560
X1116 VSS VDD 500 VDD 491 VSS sky130_fd_sc_hd__inv_8 $T=96600 204000 0 0 $X=96410 $Y=203760
X1117 VSS VDD 566 VDD 584 VSS sky130_fd_sc_hd__inv_8 $T=106260 84320 1 0 $X=106070 $Y=81360
X1118 VSS VDD 478 VDD 585 VSS sky130_fd_sc_hd__inv_8 $T=109480 122400 0 0 $X=109290 $Y=122160
X1119 VSS VDD 607 VDD 573 VSS sky130_fd_sc_hd__inv_8 $T=111780 78880 1 0 $X=111590 $Y=75920
X1120 VSS VDD SCAN_IN<16> VDD 589 VSS sky130_fd_sc_hd__inv_8 $T=117300 111520 1 0 $X=117110 $Y=108560
X1121 VSS VDD SCAN_IN<15> VDD 644 VSS sky130_fd_sc_hd__inv_8 $T=118220 116960 1 0 $X=118030 $Y=114000
X1122 VSS VDD 632 VDD 598 VSS sky130_fd_sc_hd__inv_8 $T=121900 95200 1 0 $X=121710 $Y=92240
X1123 VSS VDD 657 VDD 631 VSS sky130_fd_sc_hd__inv_8 $T=124200 29920 1 0 $X=124010 $Y=26960
X1124 VSS VDD 619 VDD 675 VSS sky130_fd_sc_hd__inv_8 $T=126500 182240 0 0 $X=126310 $Y=182000
X1125 VSS VDD SCAN_IN<14> VDD 693 VSS sky130_fd_sc_hd__inv_8 $T=133400 138720 1 0 $X=133210 $Y=135760
X1126 VSS VDD 692 VDD 706 VSS sky130_fd_sc_hd__inv_8 $T=134320 214880 0 0 $X=134130 $Y=214640
X1127 VSS VDD 713 VDD 646 VSS sky130_fd_sc_hd__inv_8 $T=136160 204000 0 0 $X=135970 $Y=203760
X1128 VSS VDD 678 VDD 680 VSS sky130_fd_sc_hd__inv_8 $T=137540 160480 1 0 $X=137350 $Y=157520
X1129 VSS VDD 673 VDD 750 VSS sky130_fd_sc_hd__inv_8 $T=138920 171360 1 0 $X=138730 $Y=168400
X1130 VSS VDD 719 VDD 700 VSS sky130_fd_sc_hd__inv_8 $T=141680 24480 1 0 $X=141490 $Y=21520
X1131 VSS VDD 736 VDD 768 VSS sky130_fd_sc_hd__inv_8 $T=143520 95200 1 0 $X=143330 $Y=92240
X1132 VSS VDD 731 VDD 520 VSS sky130_fd_sc_hd__inv_8 $T=144440 73440 1 0 $X=144250 $Y=70480
X1133 VSS VDD 677 VDD 846 VSS sky130_fd_sc_hd__inv_8 $T=162380 138720 0 0 $X=162190 $Y=138480
X1134 VSS VDD 558 VDD 798 VSS sky130_fd_sc_hd__inv_8 $T=166060 198560 0 0 $X=165870 $Y=198320
X1135 VSS VDD 532 VDD 481 VSS sky130_fd_sc_hd__inv_8 $T=170200 176800 1 0 $X=170010 $Y=173840
X1136 VSS VDD 879 VDD 815 VSS sky130_fd_sc_hd__inv_8 $T=171580 51680 1 0 $X=171390 $Y=48720
X1137 VSS VDD 893 VDD 900 VSS sky130_fd_sc_hd__inv_8 $T=175720 127840 0 0 $X=175530 $Y=127600
X1138 VSS VDD 834 VDD 873 VSS sky130_fd_sc_hd__inv_8 $T=175720 193120 1 0 $X=175530 $Y=190160
X1139 VSS VDD 863 VDD 877 VSS sky130_fd_sc_hd__inv_8 $T=176180 214880 0 0 $X=175990 $Y=214640
X1140 VSS VDD 904 VDD 749 VSS sky130_fd_sc_hd__inv_8 $T=179400 57120 0 0 $X=179210 $Y=56880
X1141 VSS VDD 823 VDD 752 VSS sky130_fd_sc_hd__inv_8 $T=180320 209440 1 0 $X=180130 $Y=206480
X1142 VSS VDD 771 VDD 784 VSS sky130_fd_sc_hd__inv_8 $T=185840 62560 0 0 $X=185650 $Y=62320
X1143 VSS VDD 956 VDD 888 VSS sky130_fd_sc_hd__inv_8 $T=190900 78880 1 0 $X=190710 $Y=75920
X1144 VSS VDD SCAN_IN<3> VDD 965 VSS sky130_fd_sc_hd__inv_8 $T=196880 204000 1 0 $X=196690 $Y=201040
X1145 VSS VDD 913 VDD 967 VSS sky130_fd_sc_hd__inv_8 $T=197800 187680 1 0 $X=197610 $Y=184720
X1146 VSS VDD 960 VDD 1033 VSS sky130_fd_sc_hd__inv_8 $T=205160 204000 1 0 $X=204970 $Y=201040
X1147 VSS VDD 940 VDD 727 VSS sky130_fd_sc_hd__inv_8 $T=205620 160480 1 0 $X=205430 $Y=157520
X1148 VSS VDD 1011 VDD 990 VSS sky130_fd_sc_hd__inv_8 $T=207920 220320 0 0 $X=207730 $Y=220080
X1149 VSS VDD 795 VDD 671 VSS sky130_fd_sc_hd__inv_8 $T=208380 225760 1 0 $X=208190 $Y=222800
X1150 VSS VDD 765 VDD 1024 VSS sky130_fd_sc_hd__inv_8 $T=209300 29920 0 0 $X=209110 $Y=29680
X1151 VSS VDD 49 84 ICV_13 $T=11960 29920 1 0 $X=11770 $Y=26960
X1152 VSS VDD 130 SCAN_IN<10> ICV_13 $T=31280 122400 1 0 $X=31090 $Y=119440
X1153 VSS VDD 186 224 ICV_13 $T=39100 57120 1 0 $X=38910 $Y=54160
X1154 VSS VDD 295 248 ICV_13 $T=49220 144160 1 0 $X=49030 $Y=141200
X1155 VSS VDD 397 430 ICV_13 $T=82340 29920 1 0 $X=82150 $Y=26960
X1156 VSS VDD 418 SCAN_IN<7> ICV_13 $T=82800 19040 1 0 $X=82610 $Y=16080
X1157 VSS VDD 326 17 ICV_13 $T=84180 106080 1 0 $X=83990 $Y=103120
X1158 VSS VDD 50 SCAN_IN<9> ICV_13 $T=91080 29920 1 0 $X=90890 $Y=26960
X1159 VSS VDD 716 702 ICV_13 $T=138000 100640 0 0 $X=137810 $Y=100400
X1160 VSS VDD 758 SCAN_IN<13> ICV_13 $T=144440 138720 1 0 $X=144250 $Y=135760
X1161 VSS VDD 464 747 ICV_13 $T=147200 220320 0 0 $X=147010 $Y=220080
X1162 VSS VDD 839 791 ICV_13 $T=166060 160480 1 0 $X=165870 $Y=157520
X1163 VSS VDD 867 881 ICV_13 $T=172040 89760 1 0 $X=171850 $Y=86800
X1164 VSS VDD 634 855 ICV_13 $T=172500 225760 1 0 $X=172310 $Y=222800
X1165 VSS VDD 909 923 ICV_13 $T=180320 116960 1 0 $X=180130 $Y=114000
X1166 VSS VDD 935 SCAN_IN<6> ICV_13 $T=180320 225760 1 0 $X=180130 $Y=222800
X1167 VSS VDD 946 801 ICV_13 $T=189980 187680 1 0 $X=189790 $Y=184720
X1168 VSS VDD 968 957 ICV_13 $T=193660 225760 1 0 $X=193470 $Y=222800
X1169 VSS VDD 422 SCAN_IN<17> ICV_13 $T=213900 95200 0 0 $X=213710 $Y=94960
X1170 VSS VDD ICV_14 $T=17020 40800 1 0 $X=16830 $Y=37840
X1171 VSS VDD ICV_14 $T=30820 204000 0 0 $X=30630 $Y=203760
X1172 VSS VDD ICV_14 $T=73140 209440 1 0 $X=72950 $Y=206480
X1173 VSS VDD ICV_14 $T=129260 62560 1 0 $X=129070 $Y=59600
X1174 VSS VDD ICV_14 $T=157320 89760 1 0 $X=157130 $Y=86800
X1175 VSS VDD ICV_14 $T=157320 106080 1 0 $X=157130 $Y=103120
X1176 VSS VDD ICV_14 $T=213440 187680 1 0 $X=213250 $Y=184720
X1177 VSS VDD ICV_14 $T=213440 204000 1 0 $X=213250 $Y=201040
X1178 VSS VDD 26 ICV_15 $T=7820 95200 1 0 $X=7630 $Y=92240
X1179 VSS VDD 11 ICV_15 $T=7820 106080 1 0 $X=7630 $Y=103120
X1180 VSS VDD 29 ICV_15 $T=7820 106080 0 0 $X=7630 $Y=105840
X1181 VSS VDD 62 ICV_15 $T=10120 57120 0 0 $X=9930 $Y=56880
X1182 VSS VDD 78 ICV_15 $T=14720 193120 1 0 $X=14530 $Y=190160
X1183 VSS VDD 65 ICV_15 $T=15640 193120 0 0 $X=15450 $Y=192880
X1184 VSS VDD 49 ICV_15 $T=16560 19040 1 0 $X=16370 $Y=16080
X1185 VSS VDD 80 ICV_15 $T=16560 46240 1 0 $X=16370 $Y=43280
X1186 VSS VDD 98 ICV_15 $T=21160 111520 0 0 $X=20970 $Y=111280
X1187 VSS VDD 113 ICV_15 $T=21160 133280 1 0 $X=20970 $Y=130320
X1188 VSS VDD 123 ICV_15 $T=21160 198560 1 0 $X=20970 $Y=195600
X1189 VSS VDD 132 ICV_15 $T=22080 182240 1 0 $X=21890 $Y=179280
X1190 VSS VDD 129 ICV_15 $T=23920 68000 0 0 $X=23730 $Y=67760
X1191 VSS VDD 119 ICV_15 $T=25300 46240 0 0 $X=25110 $Y=46000
X1192 VSS VDD 164 ICV_15 $T=27140 68000 1 0 $X=26950 $Y=65040
X1193 VSS VDD 88 ICV_15 $T=28980 35360 0 0 $X=28790 $Y=35120
X1194 VSS VDD 153 ICV_15 $T=28980 57120 0 0 $X=28790 $Y=56880
X1195 VSS VDD 173 ICV_15 $T=30820 171360 0 0 $X=30630 $Y=171120
X1196 VSS VDD 187 ICV_15 $T=34960 171360 1 0 $X=34770 $Y=168400
X1197 VSS VDD 208 ICV_15 $T=34960 209440 0 0 $X=34770 $Y=209200
X1198 VSS VDD 216 ICV_15 $T=36800 78880 1 0 $X=36610 $Y=75920
X1199 VSS VDD 241 ICV_15 $T=41860 73440 1 0 $X=41670 $Y=70480
X1200 VSS VDD 231 ICV_15 $T=42320 193120 0 0 $X=42130 $Y=192880
X1201 VSS VDD 243 ICV_15 $T=45080 62560 1 0 $X=44890 $Y=59600
X1202 VSS VDD 248 ICV_15 $T=48300 138720 0 0 $X=48110 $Y=138480
X1203 VSS VDD 317 ICV_15 $T=65320 24480 1 0 $X=65130 $Y=21520
X1204 VSS VDD 368 ICV_15 $T=65320 122400 1 0 $X=65130 $Y=119440
X1205 VSS VDD 348 ICV_15 $T=65320 182240 0 0 $X=65130 $Y=182000
X1206 VSS VDD 166 ICV_15 $T=66240 220320 1 0 $X=66050 $Y=217360
X1207 VSS VDD 382 ICV_15 $T=69920 13600 0 0 $X=69730 $Y=13360
X1208 VSS VDD 349 ICV_15 $T=70840 220320 0 0 $X=70650 $Y=220080
X1209 VSS VDD 373 ICV_15 $T=77740 46240 0 0 $X=77550 $Y=46000
X1210 VSS VDD 390 ICV_15 $T=79580 13600 0 0 $X=79390 $Y=13360
X1211 VSS VDD 281 ICV_15 $T=81420 78880 0 0 $X=81230 $Y=78640
X1212 VSS VDD 357 ICV_15 $T=81420 204000 0 0 $X=81230 $Y=203760
X1213 VSS VDD 457 ICV_15 $T=86020 187680 1 0 $X=85830 $Y=184720
X1214 VSS VDD 412 ICV_15 $T=86480 19040 0 0 $X=86290 $Y=18800
X1215 VSS VDD 455 ICV_15 $T=86480 89760 0 0 $X=86290 $Y=89520
X1216 VSS VDD 413 ICV_15 $T=86480 127840 0 0 $X=86290 $Y=127600
X1217 VSS VDD 461 ICV_15 $T=86940 122400 1 0 $X=86750 $Y=119440
X1218 VSS VDD 458 ICV_15 $T=90620 62560 1 0 $X=90430 $Y=59600
X1219 VSS VDD 431 ICV_15 $T=91080 122400 0 0 $X=90890 $Y=122160
X1220 VSS VDD 431 ICV_15 $T=94300 122400 0 0 $X=94110 $Y=122160
X1221 VSS VDD SCAN_IN<20> ICV_15 $T=96140 111520 0 0 $X=95950 $Y=111280
X1222 VSS VDD 448 ICV_15 $T=101200 116960 1 0 $X=101010 $Y=114000
X1223 VSS VDD 247 ICV_15 $T=101200 122400 1 0 $X=101010 $Y=119440
X1224 VSS VDD 509 ICV_15 $T=101660 84320 0 0 $X=101470 $Y=84080
X1225 VSS VDD 525 ICV_15 $T=103960 35360 0 0 $X=103770 $Y=35120
X1226 VSS VDD 472 ICV_15 $T=105340 127840 1 0 $X=105150 $Y=124880
X1227 VSS VDD SCAN_IN<12> ICV_15 $T=105340 138720 1 0 $X=105150 $Y=135760
X1228 VSS VDD 357 ICV_15 $T=105340 225760 1 0 $X=105150 $Y=222800
X1229 VSS VDD 562 ICV_15 $T=105800 89760 1 0 $X=105610 $Y=86800
X1230 VSS VDD 571 ICV_15 $T=107180 35360 1 0 $X=106990 $Y=32400
X1231 VSS VDD 574 ICV_15 $T=107640 68000 1 0 $X=107450 $Y=65040
X1232 VSS VDD 554 ICV_15 $T=108100 13600 0 0 $X=107910 $Y=13360
X1233 VSS VDD SCAN_IN<9> ICV_15 $T=109020 19040 0 0 $X=108830 $Y=18800
X1234 VSS VDD 522 ICV_15 $T=111320 29920 0 0 $X=111130 $Y=29680
X1235 VSS VDD SCAN_IN<12> ICV_15 $T=112700 133280 0 0 $X=112510 $Y=133040
X1236 VSS VDD 460 ICV_15 $T=112700 160480 0 0 $X=112510 $Y=160240
X1237 VSS VDD 531 ICV_15 $T=114080 122400 1 0 $X=113890 $Y=119440
X1238 VSS VDD 565 ICV_15 $T=114540 51680 0 0 $X=114350 $Y=51440
X1239 VSS VDD 605 ICV_15 $T=114540 122400 0 0 $X=114350 $Y=122160
X1240 VSS VDD 565 ICV_15 $T=115000 89760 0 0 $X=114810 $Y=89520
X1241 VSS VDD SCAN_IN<15> ICV_15 $T=119140 111520 0 0 $X=118950 $Y=111280
X1242 VSS VDD 109 ICV_15 $T=119140 144160 0 0 $X=118950 $Y=143920
X1243 VSS VDD 631 ICV_15 $T=120980 29920 1 0 $X=120790 $Y=26960
X1244 VSS VDD 632 ICV_15 $T=121900 89760 0 0 $X=121710 $Y=89520
X1245 VSS VDD 658 ICV_15 $T=123280 106080 1 0 $X=123090 $Y=103120
X1246 VSS VDD 661 ICV_15 $T=123740 111520 1 0 $X=123550 $Y=108560
X1247 VSS VDD 416 ICV_15 $T=126960 127840 1 0 $X=126770 $Y=124880
X1248 VSS VDD 641 ICV_15 $T=126960 209440 0 0 $X=126770 $Y=209200
X1249 VSS VDD 623 ICV_15 $T=128800 40800 0 0 $X=128610 $Y=40560
X1250 VSS VDD 670 ICV_15 $T=128800 68000 1 0 $X=128610 $Y=65040
X1251 VSS VDD 681 ICV_15 $T=128800 193120 1 0 $X=128610 $Y=190160
X1252 VSS VDD 682 ICV_15 $T=128800 198560 1 0 $X=128610 $Y=195600
X1253 VSS VDD 673 ICV_15 $T=131100 149600 0 0 $X=130910 $Y=149360
X1254 VSS VDD 673 ICV_15 $T=133400 155040 1 0 $X=133210 $Y=152080
X1255 VSS VDD 691 ICV_15 $T=133860 193120 0 0 $X=133670 $Y=192880
X1256 VSS VDD 706 ICV_15 $T=133860 225760 1 0 $X=133670 $Y=222800
X1257 VSS VDD 705 ICV_15 $T=136160 127840 1 0 $X=135970 $Y=124880
X1258 VSS VDD 700 ICV_15 $T=137540 19040 0 0 $X=137350 $Y=18800
X1259 VSS VDD 702 ICV_15 $T=141220 106080 0 0 $X=141030 $Y=105840
X1260 VSS VDD 719 ICV_15 $T=143060 19040 0 0 $X=142870 $Y=18800
X1261 VSS VDD 754 ICV_15 $T=143060 40800 1 0 $X=142870 $Y=37840
X1262 VSS VDD 509 ICV_15 $T=143060 73440 0 0 $X=142870 $Y=73200
X1263 VSS VDD SCAN_IN<18> ICV_15 $T=143060 78880 0 0 $X=142870 $Y=78640
X1264 VSS VDD SCAN_IN<12> ICV_15 $T=143060 138720 0 0 $X=142870 $Y=138480
X1265 VSS VDD 761 ICV_15 $T=144440 160480 1 0 $X=144250 $Y=157520
X1266 VSS VDD 676 ICV_15 $T=146280 35360 1 0 $X=146090 $Y=32400
X1267 VSS VDD 750 ICV_15 $T=146280 182240 1 0 $X=146090 $Y=179280
X1268 VSS VDD 743 ICV_15 $T=148120 122400 1 0 $X=147930 $Y=119440
X1269 VSS VDD 633 ICV_15 $T=148580 204000 1 0 $X=148390 $Y=201040
X1270 VSS VDD 731 ICV_15 $T=149500 73440 0 0 $X=149310 $Y=73200
X1271 VSS VDD SCAN_IN<16> ICV_15 $T=156400 100640 0 0 $X=156210 $Y=100400
X1272 VSS VDD 764 ICV_15 $T=157320 19040 1 0 $X=157130 $Y=16080
X1273 VSS VDD 783 ICV_15 $T=157320 149600 1 0 $X=157130 $Y=146640
X1274 VSS VDD 747 ICV_15 $T=157320 204000 0 0 $X=157130 $Y=203760
X1275 VSS VDD 783 ICV_15 $T=161460 68000 1 0 $X=161270 $Y=65040
X1276 VSS VDD 503 ICV_15 $T=161460 78880 1 0 $X=161270 $Y=75920
X1277 VSS VDD 596 ICV_15 $T=161460 116960 1 0 $X=161270 $Y=114000
X1278 VSS VDD 835 ICV_15 $T=162840 133280 1 0 $X=162650 $Y=130320
X1279 VSS VDD 798 ICV_15 $T=168820 204000 0 0 $X=168630 $Y=203760
X1280 VSS VDD 842 ICV_15 $T=169280 29920 0 0 $X=169090 $Y=29680
X1281 VSS VDD 851 ICV_15 $T=170200 133280 1 0 $X=170010 $Y=130320
X1282 VSS VDD 891 ICV_15 $T=174340 138720 1 0 $X=174150 $Y=135760
X1283 VSS VDD 895 ICV_15 $T=174340 182240 1 0 $X=174150 $Y=179280
X1284 VSS VDD 888 ICV_15 $T=176180 78880 1 0 $X=175990 $Y=75920
X1285 VSS VDD 765 ICV_15 $T=178480 57120 1 0 $X=178290 $Y=54160
X1286 VSS VDD 921 ICV_15 $T=180780 95200 1 0 $X=180590 $Y=92240
X1287 VSS VDD 893 ICV_15 $T=180780 127840 0 0 $X=180590 $Y=127600
X1288 VSS VDD 932 ICV_15 $T=182160 176800 1 0 $X=181970 $Y=173840
X1289 VSS VDD 934 ICV_15 $T=183540 100640 1 0 $X=183350 $Y=97680
X1290 VSS VDD 902 ICV_15 $T=184920 35360 1 0 $X=184730 $Y=32400
X1291 VSS VDD 759 ICV_15 $T=184920 149600 1 0 $X=184730 $Y=146640
X1292 VSS VDD 864 ICV_15 $T=185380 19040 1 0 $X=185190 $Y=16080
X1293 VSS VDD 848 ICV_15 $T=189520 95200 1 0 $X=189330 $Y=92240
X1294 VSS VDD 712 ICV_15 $T=190440 122400 0 0 $X=190250 $Y=122160
X1295 VSS VDD 892 ICV_15 $T=190440 127840 1 0 $X=190250 $Y=124880
X1296 VSS VDD 956 ICV_15 $T=191360 73440 0 0 $X=191170 $Y=73200
X1297 VSS VDD 774 ICV_15 $T=192280 95200 0 0 $X=192090 $Y=94960
X1298 VSS VDD 915 ICV_15 $T=192280 144160 0 0 $X=192090 $Y=143920
X1299 VSS VDD 976 ICV_15 $T=195500 95200 0 0 $X=195310 $Y=94960
X1300 VSS VDD 727 ICV_15 $T=195960 149600 0 0 $X=195770 $Y=149360
X1301 VSS VDD 912 ICV_15 $T=197340 57120 0 0 $X=197150 $Y=56880
X1302 VSS VDD 969 ICV_15 $T=198720 29920 0 0 $X=198530 $Y=29680
X1303 VSS VDD 723 ICV_15 $T=199180 149600 0 0 $X=198990 $Y=149360
X1304 VSS VDD SCAN_IN<0> ICV_15 $T=199180 155040 0 0 $X=198990 $Y=154800
X1305 VSS VDD 992 ICV_15 $T=201940 204000 1 0 $X=201750 $Y=201040
X1306 VSS VDD 972 ICV_15 $T=202860 127840 1 0 $X=202670 $Y=124880
X1307 VSS VDD 986 ICV_15 $T=203320 84320 0 0 $X=203130 $Y=84080
X1308 VSS VDD 913 ICV_15 $T=203320 193120 0 0 $X=203130 $Y=192880
X1309 VSS VDD 701 ICV_15 $T=204240 51680 1 0 $X=204050 $Y=48720
X1310 VSS VDD 1024 ICV_15 $T=207000 24480 0 0 $X=206810 $Y=24240
X1311 VSS VDD 1010 ICV_15 $T=207920 209440 0 0 $X=207730 $Y=209200
X1312 VSS VDD 1037 ICV_15 $T=212980 40800 1 0 $X=212790 $Y=37840
X1313 VSS VDD 1038 ICV_15 $T=212980 62560 1 0 $X=212790 $Y=59600
X1314 VSS VDD 988 ICV_15 $T=212980 116960 1 0 $X=212790 $Y=114000
X1315 VSS VDD 163 ICV_16 $T=30820 29920 0 0 $X=30630 $Y=29680
X1316 VSS VDD 19 ICV_16 $T=30820 40800 0 0 $X=30630 $Y=40560
X1317 VSS VDD 57 ICV_16 $T=30820 149600 0 0 $X=30630 $Y=149360
X1318 VSS VDD 132 ICV_16 $T=30820 182240 0 0 $X=30630 $Y=182000
X1319 VSS VDD 260 ICV_16 $T=45080 35360 1 0 $X=44890 $Y=32400
X1320 VSS VDD 236 ICV_16 $T=45080 68000 1 0 $X=44890 $Y=65040
X1321 VSS VDD 263 ICV_16 $T=45080 160480 1 0 $X=44890 $Y=157520
X1322 VSS VDD 84 ICV_16 $T=58880 24480 0 0 $X=58690 $Y=24240
X1323 VSS VDD 310 ICV_16 $T=58880 220320 0 0 $X=58690 $Y=220080
X1324 VSS VDD 412 ICV_16 $T=86940 24480 0 0 $X=86750 $Y=24240
X1325 VSS VDD 441 ICV_16 $T=86940 176800 0 0 $X=86750 $Y=176560
X1326 VSS VDD 529 ICV_16 $T=101200 51680 1 0 $X=101010 $Y=48720
X1327 VSS VDD 685 ICV_16 $T=129260 182240 1 0 $X=129070 $Y=179280
X1328 VSS VDD 719 ICV_16 $T=143060 29920 0 0 $X=142870 $Y=29680
X1329 VSS VDD 807 ICV_16 $T=157320 24480 1 0 $X=157130 $Y=21520
X1330 VSS VDD 797 ICV_16 $T=157320 46240 1 0 $X=157130 $Y=43280
X1331 VSS VDD 785 ICV_16 $T=157320 155040 1 0 $X=157130 $Y=152080
X1332 VSS VDD 905 ICV_16 $T=185380 176800 1 0 $X=185190 $Y=173840
X1333 VSS VDD SCAN_IN<5> ICV_16 $T=199180 78880 0 0 $X=198990 $Y=78640
X1334 VSS VDD 987 ICV_16 $T=199180 100640 0 0 $X=198990 $Y=100400
X1335 VSS VDD 723 ICV_16 $T=199180 133280 0 0 $X=198990 $Y=133040
X1336 VSS VDD 819 ICV_16 $T=199180 144160 0 0 $X=198990 $Y=143920
X1337 VSS VDD 904 ICV_16 $T=202400 13600 1 0 $X=202210 $Y=10640
X1338 VSS VDD 1051 ICV_16 $T=213440 24480 1 0 $X=213250 $Y=21520
X1339 VSS VDD 1035 ICV_16 $T=213440 122400 1 0 $X=213250 $Y=119440
X1340 VSS VDD 1042 ICV_16 $T=213440 155040 1 0 $X=213250 $Y=152080
X1341 VSS VDD ICV_17 $T=11960 171360 0 0 $X=11770 $Y=171120
X1342 VSS VDD ICV_17 $T=24380 225760 1 0 $X=24190 $Y=222800
X1343 VSS VDD ICV_17 $T=25300 57120 1 0 $X=25110 $Y=54160
X1344 VSS VDD ICV_17 $T=37720 165920 1 0 $X=37530 $Y=162960
X1345 VSS VDD ICV_17 $T=39100 198560 1 0 $X=38910 $Y=195600
X1346 VSS VDD ICV_17 $T=40940 171360 0 0 $X=40750 $Y=171120
X1347 VSS VDD ICV_17 $T=41860 214880 0 0 $X=41670 $Y=214640
X1348 VSS VDD ICV_17 $T=68080 144160 0 0 $X=67890 $Y=143920
X1349 VSS VDD ICV_17 $T=78660 225760 1 0 $X=78470 $Y=222800
X1350 VSS VDD ICV_17 $T=80960 138720 0 0 $X=80770 $Y=138480
X1351 VSS VDD ICV_17 $T=93840 182240 0 0 $X=93650 $Y=182000
X1352 VSS VDD ICV_17 $T=106720 171360 1 0 $X=106530 $Y=168400
X1353 VSS VDD ICV_17 $T=123740 73440 1 0 $X=123550 $Y=70480
X1354 VSS VDD ICV_17 $T=143060 68000 1 0 $X=142870 $Y=65040
X1355 VSS VDD ICV_17 $T=179860 193120 1 0 $X=179670 $Y=190160
X1356 VSS VDD ICV_17 $T=179860 204000 1 0 $X=179670 $Y=201040
X1357 VSS VDD ICV_17 $T=180320 214880 0 0 $X=180130 $Y=214640
X1358 VSS VDD ICV_17 $T=192740 89760 1 0 $X=192550 $Y=86800
X1359 VSS VDD ICV_17 $T=193660 214880 1 0 $X=193470 $Y=211920
X1360 VSS VDD ICV_17 $T=207460 106080 1 0 $X=207270 $Y=103120
X1361 VSS VDD ICV_17 $T=213440 29920 0 0 $X=213250 $Y=29680
X1362 VSS VDD ICV_18 $T=16100 51680 1 0 $X=15910 $Y=48720
X1363 VSS VDD ICV_18 $T=16100 73440 1 0 $X=15910 $Y=70480
X1364 VSS VDD ICV_18 $T=16100 160480 1 0 $X=15910 $Y=157520
X1365 VSS VDD ICV_18 $T=44160 111520 1 0 $X=43970 $Y=108560
X1366 VSS VDD ICV_18 $T=44160 138720 1 0 $X=43970 $Y=135760
X1367 VSS VDD ICV_18 $T=44160 144160 1 0 $X=43970 $Y=141200
X1368 VSS VDD ICV_18 $T=44160 187680 1 0 $X=43970 $Y=184720
X1369 VSS VDD ICV_18 $T=72220 24480 1 0 $X=72030 $Y=21520
X1370 VSS VDD ICV_18 $T=72220 51680 1 0 $X=72030 $Y=48720
X1371 VSS VDD ICV_18 $T=72220 73440 1 0 $X=72030 $Y=70480
X1372 VSS VDD ICV_18 $T=72220 106080 1 0 $X=72030 $Y=103120
X1373 VSS VDD ICV_18 $T=72220 122400 1 0 $X=72030 $Y=119440
X1374 VSS VDD ICV_18 $T=72220 144160 1 0 $X=72030 $Y=141200
X1375 VSS VDD ICV_18 $T=100280 40800 1 0 $X=100090 $Y=37840
X1376 VSS VDD ICV_18 $T=100280 89760 1 0 $X=100090 $Y=86800
X1377 VSS VDD ICV_18 $T=128340 40800 1 0 $X=128150 $Y=37840
X1378 VSS VDD ICV_18 $T=128340 46240 1 0 $X=128150 $Y=43280
X1379 VSS VDD ICV_18 $T=128340 100640 1 0 $X=128150 $Y=97680
X1380 VSS VDD ICV_18 $T=156400 35360 1 0 $X=156210 $Y=32400
X1381 VSS VDD ICV_18 $T=156400 138720 1 0 $X=156210 $Y=135760
X1382 VSS VDD ICV_18 $T=156400 209440 1 0 $X=156210 $Y=206480
X1383 VSS VDD ICV_18 $T=156400 220320 1 0 $X=156210 $Y=217360
X1384 VSS VDD ICV_18 $T=170200 198560 0 0 $X=170010 $Y=198320
X1385 VSS VDD ICV_18 $T=184460 73440 1 0 $X=184270 $Y=70480
X1386 VSS VDD ICV_18 $T=184460 160480 1 0 $X=184270 $Y=157520
X1387 VSS VDD ICV_18 $T=184460 171360 1 0 $X=184270 $Y=168400
X1388 VSS VDD ICV_18 $T=184460 187680 1 0 $X=184270 $Y=184720
X1389 VSS VDD ICV_18 $T=201480 225760 0 0 $X=201290 $Y=225520
X1390 VSS VDD ICV_19 $T=212520 19040 1 0 $X=212330 $Y=16080
X1391 VSS VDD ICV_19 $T=212520 51680 1 0 $X=212330 $Y=48720
X1392 VSS VDD ICV_19 $T=212520 73440 1 0 $X=212330 $Y=70480
X1393 VSS VDD ICV_19 $T=212520 78880 1 0 $X=212330 $Y=75920
X1394 VSS VDD ICV_19 $T=212520 100640 1 0 $X=212330 $Y=97680
X1395 VSS VDD ICV_19 $T=212520 138720 1 0 $X=212330 $Y=135760
X1396 VSS VDD ICV_19 $T=212520 176800 1 0 $X=212330 $Y=173840
X1397 VSS VDD ICV_19 $T=212520 193120 1 0 $X=212330 $Y=190160
X1398 VSS VDD ICV_19 $T=212520 225760 1 0 $X=212330 $Y=222800
X1399 VSS VDD 38 ICV_20 $T=12420 19040 1 0 $X=12230 $Y=16080
X1400 VSS VDD 55 ICV_20 $T=15640 84320 1 0 $X=15450 $Y=81360
X1401 VSS VDD 26 ICV_20 $T=15640 84320 0 0 $X=15450 $Y=84080
X1402 VSS VDD 25 ICV_20 $T=15640 106080 1 0 $X=15450 $Y=103120
X1403 VSS VDD 10 ICV_20 $T=16100 68000 1 0 $X=15910 $Y=65040
X1404 VSS VDD 91 ICV_20 $T=19320 100640 0 0 $X=19130 $Y=100400
X1405 VSS VDD 61 ICV_20 $T=29440 24480 0 0 $X=29250 $Y=24240
X1406 VSS VDD 159 ICV_20 $T=32200 116960 1 0 $X=32010 $Y=114000
X1407 VSS VDD 162 ICV_20 $T=39100 220320 0 0 $X=38910 $Y=220080
X1408 VSS VDD 64 ICV_20 $T=40020 100640 1 0 $X=39830 $Y=97680
X1409 VSS VDD 255 ICV_20 $T=43700 95200 1 0 $X=43510 $Y=92240
X1410 VSS VDD 217 ICV_20 $T=43700 100640 1 0 $X=43510 $Y=97680
X1411 VSS VDD 214 ICV_20 $T=43700 106080 1 0 $X=43510 $Y=103120
X1412 VSS VDD 229 ICV_20 $T=44160 84320 1 0 $X=43970 $Y=81360
X1413 VSS VDD 222 ICV_20 $T=45080 176800 0 0 $X=44890 $Y=176560
X1414 VSS VDD 17 ICV_20 $T=55660 111520 0 0 $X=55470 $Y=111280
X1415 VSS VDD 297 ICV_20 $T=56580 220320 1 0 $X=56390 $Y=217360
X1416 VSS VDD 291 ICV_20 $T=57960 198560 1 0 $X=57770 $Y=195600
X1417 VSS VDD 341 ICV_20 $T=66700 78880 0 0 $X=66510 $Y=78640
X1418 VSS VDD 388 ICV_20 $T=70380 133280 1 0 $X=70190 $Y=130320
X1419 VSS VDD 397 ICV_20 $T=71760 29920 1 0 $X=71570 $Y=26960
X1420 VSS VDD 376 ICV_20 $T=72220 19040 1 0 $X=72030 $Y=16080
X1421 VSS VDD 353 ICV_20 $T=72220 176800 1 0 $X=72030 $Y=173840
X1422 VSS VDD 135 ICV_20 $T=74980 127840 0 0 $X=74790 $Y=127600
X1423 VSS VDD 425 ICV_20 $T=81880 155040 0 0 $X=81690 $Y=154800
X1424 VSS VDD 471 ICV_20 $T=88320 144160 1 0 $X=88130 $Y=141200
X1425 VSS VDD 468 ICV_20 $T=90160 155040 1 0 $X=89970 $Y=152080
X1426 VSS VDD 415 ICV_20 $T=95220 78880 1 0 $X=95030 $Y=75920
X1427 VSS VDD 512 ICV_20 $T=115460 171360 1 0 $X=115270 $Y=168400
X1428 VSS VDD 561 ICV_20 $T=120060 144160 1 0 $X=119870 $Y=141200
X1429 VSS VDD 600 ICV_20 $T=120980 165920 1 0 $X=120790 $Y=162960
X1430 VSS VDD 628 ICV_20 $T=128340 51680 1 0 $X=128150 $Y=48720
X1431 VSS VDD 663 ICV_20 $T=128340 225760 1 0 $X=128150 $Y=222800
X1432 VSS VDD 678 ICV_20 $T=136160 160480 0 0 $X=135970 $Y=160240
X1433 VSS VDD 739 ICV_20 $T=139840 127840 0 0 $X=139650 $Y=127600
X1434 VSS VDD 578 ICV_20 $T=142600 57120 1 0 $X=142410 $Y=54160
X1435 VSS VDD 677 ICV_20 $T=155020 111520 0 0 $X=154830 $Y=111280
X1436 VSS VDD 799 ICV_20 $T=156400 144160 1 0 $X=156210 $Y=141200
X1437 VSS VDD 786 ICV_20 $T=163760 209440 1 0 $X=163570 $Y=206480
X1438 VSS VDD 791 ICV_20 $T=166060 155040 0 0 $X=165870 $Y=154800
X1439 VSS VDD 855 ICV_20 $T=166520 220320 1 0 $X=166330 $Y=217360
X1440 VSS VDD 840 ICV_20 $T=170660 182240 1 0 $X=170470 $Y=179280
X1441 VSS VDD 17 ICV_20 $T=177560 155040 0 0 $X=177370 $Y=154800
X1442 VSS VDD 833 ICV_20 $T=179860 100640 1 0 $X=179670 $Y=97680
X1443 VSS VDD 851 ICV_20 $T=181240 133280 0 0 $X=181050 $Y=133040
X1444 VSS VDD SCAN_IN<5> ICV_20 $T=195960 171360 0 0 $X=195770 $Y=171120
X1445 VSS VDD 937 ICV_20 $T=196420 35360 0 0 $X=196230 $Y=35120
X1446 VSS VDD 956 ICV_20 $T=196420 73440 0 0 $X=196230 $Y=73200
X1447 VSS VDD 981 ICV_20 $T=197800 13600 0 0 $X=197610 $Y=13360
X1448 VSS VDD 913 ICV_20 $T=197800 182240 0 0 $X=197610 $Y=182000
X1449 VSS VDD 1015 ICV_20 $T=207000 62560 0 0 $X=206810 $Y=62320
X1450 VSS VDD 1045 ICV_20 $T=212060 29920 1 0 $X=211870 $Y=26960
X1451 VSS VDD 1023 ICV_20 $T=212060 198560 1 0 $X=211870 $Y=195600
X1452 VSS VDD 671 ICV_20 $T=212060 220320 1 0 $X=211870 $Y=217360
X1453 VSS VDD 1035 ICV_20 $T=212520 133280 1 0 $X=212330 $Y=130320
X1454 VSS 21 10 ICV_21 $T=7820 35360 1 0 $X=7630 $Y=32400
X1455 VSS 37 29 ICV_21 $T=8280 89760 1 0 $X=8090 $Y=86800
X1456 VSS 43 20 ICV_21 $T=8740 68000 0 0 $X=8550 $Y=67760
X1457 VSS 49 70 ICV_21 $T=9200 13600 1 0 $X=9010 $Y=10640
X1458 VSS 85 61 ICV_21 $T=14260 40800 1 0 $X=14070 $Y=37840
X1459 VSS 72 49 ICV_21 $T=15180 24480 1 0 $X=14990 $Y=21520
X1460 VSS 90 95 ICV_21 $T=15180 165920 0 0 $X=14990 $Y=165680
X1461 VSS 89 20 ICV_21 $T=15640 78880 0 0 $X=15450 $Y=78640
X1462 VSS 93 109 ICV_21 $T=16560 133280 0 0 $X=16370 $Y=133040
X1463 VSS 97 111 ICV_21 $T=17020 198560 0 0 $X=16830 $Y=198320
X1464 VSS 107 80 ICV_21 $T=18400 51680 0 0 $X=18210 $Y=51440
X1465 VSS 61 128 ICV_21 $T=20240 35360 0 0 $X=20050 $Y=35120
X1466 VSS 102 90 ICV_21 $T=20240 171360 0 0 $X=20050 $Y=171120
X1467 VSS 110 101 ICV_21 $T=20240 220320 0 0 $X=20050 $Y=220080
X1468 VSS 61 85 ICV_21 $T=21160 40800 0 0 $X=20970 $Y=40560
X1469 VSS 108 107 ICV_21 $T=21160 62560 0 0 $X=20970 $Y=62320
X1470 VSS 151 145 ICV_21 $T=26220 214880 1 0 $X=26030 $Y=211920
X1471 VSS 152 120 ICV_21 $T=27600 100640 0 0 $X=27410 $Y=100400
X1472 VSS 65 145 ICV_21 $T=28060 204000 0 0 $X=27870 $Y=203760
X1473 VSS 177 152 ICV_21 $T=28520 106080 0 0 $X=28330 $Y=105840
X1474 VSS 87 143 ICV_21 $T=28980 182240 1 0 $X=28790 $Y=179280
X1475 VSS 146 127 ICV_21 $T=29900 214880 0 0 $X=29710 $Y=214640
X1476 VSS 183 16 ICV_21 $T=29900 220320 0 0 $X=29710 $Y=220080
X1477 VSS 186 192 ICV_21 $T=31280 62560 1 0 $X=31090 $Y=59600
X1478 VSS 187 188 ICV_21 $T=31280 149600 1 0 $X=31090 $Y=146640
X1479 VSS 165 201 ICV_21 $T=31740 89760 1 0 $X=31550 $Y=86800
X1480 VSS 140 91 ICV_21 $T=32200 100640 1 0 $X=32010 $Y=97680
X1481 VSS 191 20 ICV_21 $T=34960 13600 0 0 $X=34770 $Y=13360
X1482 VSS 148 219 ICV_21 $T=34960 149600 0 0 $X=34770 $Y=149360
X1483 VSS 156 221 ICV_21 $T=35420 133280 1 0 $X=35230 $Y=130320
X1484 VSS 194 226 ICV_21 $T=36340 111520 0 0 $X=36150 $Y=111280
X1485 VSS 222 173 ICV_21 $T=38180 171360 0 0 $X=37990 $Y=171120
X1486 VSS 184 138 ICV_21 $T=39100 214880 0 0 $X=38910 $Y=214640
X1487 VSS 232 238 ICV_21 $T=39560 29920 0 0 $X=39370 $Y=29680
X1488 VSS 161 206 ICV_21 $T=39560 187680 0 0 $X=39370 $Y=187440
X1489 VSS 250 191 ICV_21 $T=43240 29920 1 0 $X=43050 $Y=26960
X1490 VSS 252 258 ICV_21 $T=43240 155040 1 0 $X=43050 $Y=152080
X1491 VSS 253 271 ICV_21 $T=45080 149600 0 0 $X=44890 $Y=149360
X1492 VSS 161 272 ICV_21 $T=45080 198560 0 0 $X=44890 $Y=198320
X1493 VSS 271 249 ICV_21 $T=46460 182240 0 0 $X=46270 $Y=182000
X1494 VSS 225 272 ICV_21 $T=46460 209440 0 0 $X=46270 $Y=209200
X1495 VSS 274 287 ICV_21 $T=47840 24480 0 0 $X=47650 $Y=24240
X1496 VSS 284 243 ICV_21 $T=49220 68000 0 0 $X=49030 $Y=67760
X1497 VSS 119 119 ICV_21 $T=54740 73440 1 0 $X=54550 $Y=70480
X1498 VSS 250 322 ICV_21 $T=56580 35360 0 0 $X=56390 $Y=35120
X1499 VSS 275 284 ICV_21 $T=56580 62560 0 0 $X=56390 $Y=62320
X1500 VSS 295 304 ICV_21 $T=56580 133280 0 0 $X=56390 $Y=133040
X1501 VSS 325 324 ICV_21 $T=57500 160480 0 0 $X=57310 $Y=160240
X1502 VSS 310 106 ICV_21 $T=57500 204000 0 0 $X=57310 $Y=203760
X1503 VSS 327 271 ICV_21 $T=57960 149600 0 0 $X=57770 $Y=149360
X1504 VSS 310 338 ICV_21 $T=57960 176800 0 0 $X=57770 $Y=176560
X1505 VSS 150 190 ICV_21 $T=62100 198560 1 0 $X=61910 $Y=195600
X1506 VSS 168 373 ICV_21 $T=65320 62560 0 0 $X=65130 $Y=62320
X1507 VSS 107 323 ICV_21 $T=65320 73440 1 0 $X=65130 $Y=70480
X1508 VSS 367 346 ICV_21 $T=65320 106080 0 0 $X=65130 $Y=105840
X1509 VSS 327 315 ICV_21 $T=65320 144160 0 0 $X=65130 $Y=143920
X1510 VSS 339 310 ICV_21 $T=65320 187680 0 0 $X=65130 $Y=187440
X1511 VSS 348 356 ICV_21 $T=67160 149600 0 0 $X=66970 $Y=149360
X1512 VSS 238 386 ICV_21 $T=68080 24480 0 0 $X=67890 $Y=24240
X1513 VSS 245 398 ICV_21 $T=70380 209440 1 0 $X=70190 $Y=206480
X1514 VSS 391 383 ICV_21 $T=70840 29920 0 0 $X=70650 $Y=29680
X1515 VSS 125 393 ICV_21 $T=70840 78880 0 0 $X=70650 $Y=78640
X1516 VSS 394 349 ICV_21 $T=71300 187680 1 0 $X=71110 $Y=184720
X1517 VSS 275 375 ICV_21 $T=73140 68000 0 0 $X=72950 $Y=67760
X1518 VSS 407 356 ICV_21 $T=74520 160480 0 0 $X=74330 $Y=160240
X1519 VSS 338 433 ICV_21 $T=77280 176800 0 0 $X=77090 $Y=176560
X1520 VSS 388 438 ICV_21 $T=78660 122400 0 0 $X=78470 $Y=122160
X1521 VSS 416 454 ICV_21 $T=84180 78880 1 0 $X=83990 $Y=75920
X1522 VSS 373 379 ICV_21 $T=84640 46240 0 0 $X=84450 $Y=46000
X1523 VSS 448 248 ICV_21 $T=86020 144160 0 0 $X=85830 $Y=143920
X1524 VSS 475 473 ICV_21 $T=90160 133280 1 0 $X=89970 $Y=130320
X1525 VSS 337 189 ICV_21 $T=91080 182240 0 0 $X=90890 $Y=182000
X1526 VSS 484 466 ICV_21 $T=92000 95200 0 0 $X=91810 $Y=94960
X1527 VSS 489 510 ICV_21 $T=94300 51680 0 0 $X=94110 $Y=51440
X1528 VSS 486 486 ICV_21 $T=96600 144160 0 0 $X=96410 $Y=143920
X1529 VSS 516 522 ICV_21 $T=97980 19040 0 0 $X=97790 $Y=18800
X1530 VSS 519 502 ICV_21 $T=98900 46240 1 0 $X=98710 $Y=43280
X1531 VSS 436 531 ICV_21 $T=99360 127840 1 0 $X=99170 $Y=124880
X1532 VSS 526 473 ICV_21 $T=100280 144160 1 0 $X=100090 $Y=141200
X1533 VSS 466 109 ICV_21 $T=100280 149600 0 0 $X=100090 $Y=149360
X1534 VSS 535 547 ICV_21 $T=101660 204000 0 0 $X=101470 $Y=203760
X1535 VSS 532 476 ICV_21 $T=105340 165920 0 0 $X=105150 $Y=165680
X1536 VSS 513 574 ICV_21 $T=107180 40800 0 0 $X=106990 $Y=40560
X1537 VSS 573 SCAN_IN<21> ICV_21 $T=107180 100640 0 0 $X=106990 $Y=100400
X1538 VSS 577 584 ICV_21 $T=108100 78880 1 0 $X=107910 $Y=75920
X1539 VSS 596 529 ICV_21 $T=111320 62560 1 0 $X=111130 $Y=59600
X1540 VSS 570 577 ICV_21 $T=111780 51680 1 0 $X=111590 $Y=48720
X1541 VSS 337 590 ICV_21 $T=113620 171360 0 0 $X=113430 $Y=171120
X1542 VSS 618 644 ICV_21 $T=119140 116960 0 0 $X=118950 $Y=116720
X1543 VSS 634 647 ICV_21 $T=119140 220320 0 0 $X=118950 $Y=220080
X1544 VSS 640 651 ICV_21 $T=120060 176800 0 0 $X=119870 $Y=176560
X1545 VSS SCAN_IN<19> 637 ICV_21 $T=120520 68000 0 0 $X=120330 $Y=67760
X1546 VSS 641 653 ICV_21 $T=120520 187680 0 0 $X=120330 $Y=187440
X1547 VSS SCAN_IN<14> 624 ICV_21 $T=123280 127840 0 0 $X=123090 $Y=127600
X1548 VSS 534 632 ICV_21 $T=125580 46240 1 0 $X=125390 $Y=43280
X1549 VSS 548 20 ICV_21 $T=126500 78880 0 0 $X=126310 $Y=78640
X1550 VSS 534 687 ICV_21 $T=128340 57120 1 0 $X=128150 $Y=54160
X1551 VSS SCAN_IN<14> SCAN_IN<12> ICV_21 $T=131100 133280 0 0 $X=130910 $Y=133040
X1552 VSS 691 665 ICV_21 $T=135700 187680 1 0 $X=135510 $Y=184720
X1553 VSS 717 729 ICV_21 $T=142140 111520 0 0 $X=141950 $Y=111280
X1554 VSS 750 590 ICV_21 $T=142140 171360 0 0 $X=141950 $Y=171120
X1555 VSS 752 728 ICV_21 $T=142140 198560 0 0 $X=141950 $Y=198320
X1556 VSS 628 443 ICV_21 $T=147200 51680 0 0 $X=147010 $Y=51440
X1557 VSS 785 791 ICV_21 $T=150420 149600 0 0 $X=150230 $Y=149360
X1558 VSS 789 788 ICV_21 $T=152260 24480 0 0 $X=152070 $Y=24240
X1559 VSS 20 16 ICV_21 $T=155020 220320 0 0 $X=154830 $Y=220080
X1560 VSS 804 337 ICV_21 $T=156400 171360 0 0 $X=156210 $Y=171120
X1561 VSS 810 700 ICV_21 $T=159160 35360 0 0 $X=158970 $Y=35120
X1562 VSS 816 822 ICV_21 $T=159160 127840 0 0 $X=158970 $Y=127600
X1563 VSS 774 730 ICV_21 $T=161460 106080 1 0 $X=161270 $Y=103120
X1564 VSS 677 677 ICV_21 $T=161460 138720 1 0 $X=161270 $Y=135760
X1565 VSS 823 696 ICV_21 $T=163760 204000 1 0 $X=163570 $Y=201040
X1566 VSS 874 869 ICV_21 $T=169280 40800 1 0 $X=169090 $Y=37840
X1567 VSS 879 887 ICV_21 $T=170200 46240 0 0 $X=170010 $Y=46000
X1568 VSS 881 888 ICV_21 $T=170200 84320 0 0 $X=170010 $Y=84080
X1569 VSS 882 20 ICV_21 $T=170200 155040 0 0 $X=170010 $Y=154800
X1570 VSS 872 872 ICV_21 $T=170200 165920 0 0 $X=170010 $Y=165680
X1571 VSS 884 897 ICV_21 $T=170660 35360 1 0 $X=170470 $Y=32400
X1572 VSS 902 887 ICV_21 $T=175260 40800 0 0 $X=175070 $Y=40560
X1573 VSS 855 SCAN_IN<1> ICV_21 $T=175260 220320 0 0 $X=175070 $Y=220080
X1574 VSS 912 867 ICV_21 $T=177560 68000 0 0 $X=177370 $Y=67760
X1575 VSS 17 854 ICV_21 $T=177560 198560 1 0 $X=177370 $Y=195600
X1576 VSS 870 17 ICV_21 $T=178480 160480 0 0 $X=178290 $Y=160240
X1577 VSS 916 481 ICV_21 $T=178480 171360 0 0 $X=178290 $Y=171120
X1578 VSS 926 912 ICV_21 $T=181700 73440 1 0 $X=181510 $Y=70480
X1579 VSS 936 776 ICV_21 $T=184000 127840 1 0 $X=183810 $Y=124880
X1580 VSS 801 SCAN_IN<5> ICV_21 $T=184920 165920 0 0 $X=184730 $Y=165680
X1581 VSS 875 930 ICV_21 $T=188600 29920 0 0 $X=188410 $Y=29680
X1582 VSS 919 927 ICV_21 $T=188600 84320 0 0 $X=188410 $Y=84080
X1583 VSS 927 SCAN_IN<5> ICV_21 $T=189520 78880 0 0 $X=189330 $Y=78640
X1584 VSS 661 928 ICV_21 $T=192280 144160 1 0 $X=192090 $Y=141200
X1585 VSS SCAN_IN<0> 929 ICV_21 $T=193660 160480 0 0 $X=193470 $Y=160240
X1586 VSS 956 956 ICV_21 $T=195960 78880 1 0 $X=195770 $Y=75920
X1587 VSS 993 650 ICV_21 $T=198260 40800 0 0 $X=198070 $Y=40560
X1588 VSS 902 1000 ICV_21 $T=198260 51680 0 0 $X=198070 $Y=51440
X1589 VSS 1009 970 ICV_21 $T=202860 84320 1 0 $X=202670 $Y=81360
X1590 VSS 978 940 ICV_21 $T=203320 171360 0 0 $X=203130 $Y=171120
X1591 VSS 1011 795 ICV_21 $T=204240 220320 0 0 $X=204050 $Y=220080
X1592 VSS 1023 1026 ICV_21 $T=207000 182240 0 0 $X=206810 $Y=182000
X1593 VSS 1032 988 ICV_21 $T=207920 155040 0 0 $X=207730 $Y=154800
X1594 VSS 784 1041 ICV_21 $T=208380 57120 0 0 $X=208190 $Y=56880
X1595 VSS 1025 1003 ICV_21 $T=208380 160480 0 0 $X=208190 $Y=160240
X1596 VSS 984 1012 ICV_21 $T=208380 171360 1 0 $X=208190 $Y=168400
X1597 VSS 911 1037 ICV_21 $T=209300 46240 1 0 $X=209110 $Y=43280
X1598 VSS 1015 1034 ICV_21 $T=209300 68000 0 0 $X=209110 $Y=67760
X1599 VSS 1043 1049 ICV_21 $T=212060 149600 1 0 $X=211870 $Y=146640
X1600 VSS 1048 1025 ICV_21 $T=212060 165920 1 0 $X=211870 $Y=162960
X1601 VSS VDD RESET_N 38 ICV_22 $T=7820 133280 0 0 $X=7630 $Y=133040
X1602 VSS VDD 16 51 ICV_22 $T=7820 182240 1 0 $X=7630 $Y=179280
X1603 VSS VDD BB_IN 31 ICV_22 $T=10120 127840 1 0 $X=9930 $Y=124880
X1604 VSS VDD RESET_N 41 ICV_22 $T=10120 220320 1 0 $X=9930 $Y=217360
X1605 VSS VDD 227 124 ICV_22 $T=38640 13600 1 0 $X=38450 $Y=10640
X1606 VSS VDD 188 256 ICV_22 $T=48760 160480 0 0 $X=48570 $Y=160240
X1607 VSS VDD 127 258 ICV_22 $T=49220 193120 0 0 $X=49030 $Y=192880
X1608 VSS VDD 372 350 ICV_22 $T=68540 40800 0 0 $X=68350 $Y=40560
X1609 VSS VDD 345 7 ICV_22 $T=76360 95200 0 0 $X=76170 $Y=94960
X1610 VSS VDD 538 499 ICV_22 $T=104420 171360 0 0 $X=104230 $Y=171120
X1611 VSS VDD 452 520 ICV_22 $T=105340 46240 0 0 $X=105150 $Y=46000
X1612 VSS VDD 561 568 ICV_22 $T=105340 144160 0 0 $X=105150 $Y=143920
X1613 VSS VDD 623 655 ICV_22 $T=121900 19040 1 0 $X=121710 $Y=16080
X1614 VSS VDD 662 456 ICV_22 $T=123740 144160 1 0 $X=123550 $Y=141200
X1615 VSS VDD 641 690 ICV_22 $T=136160 209440 0 0 $X=135970 $Y=209200
X1616 VSS VDD 713 690 ICV_22 $T=137080 193120 0 0 $X=136890 $Y=192880
X1617 VSS VDD 765 422 ICV_22 $T=146280 89760 1 0 $X=146090 $Y=86800
X1618 VSS VDD 520 521 ICV_22 $T=150880 51680 1 0 $X=150690 $Y=48720
X1619 VSS VDD 620 862 ICV_22 $T=165600 187680 0 0 $X=165410 $Y=187440
X1620 VSS VDD 519 884 ICV_22 $T=178940 46240 1 0 $X=178750 $Y=43280
X1621 VSS VDD 1018 844 ICV_22 $T=206080 35360 1 0 $X=205890 $Y=32400
X1622 VSS VDD 976 1019 ICV_22 $T=207460 95200 1 0 $X=207270 $Y=92240
X1623 VSS VDD 1024 1036 ICV_22 $T=212520 19040 0 0 $X=212330 $Y=18800
X1624 VSS VDD ICV_23 $T=10580 35360 1 0 $X=10390 $Y=32400
X1625 VSS VDD ICV_23 $T=37720 220320 1 0 $X=37530 $Y=217360
X1626 VSS VDD ICV_23 $T=38180 133280 1 0 $X=37990 $Y=130320
X1627 VSS VDD ICV_23 $T=45080 40800 0 0 $X=44890 $Y=40560
X1628 VSS VDD ICV_23 $T=58420 40800 1 0 $X=58230 $Y=37840
X1629 VSS VDD ICV_23 $T=60720 209440 1 0 $X=60530 $Y=206480
X1630 VSS VDD ICV_23 $T=61640 187680 1 0 $X=61450 $Y=184720
X1631 VSS VDD ICV_23 $T=66700 165920 1 0 $X=66510 $Y=162960
X1632 VSS VDD ICV_23 $T=76360 198560 1 0 $X=76170 $Y=195600
X1633 VSS VDD ICV_23 $T=83720 89760 1 0 $X=83530 $Y=86800
X1634 VSS VDD ICV_23 $T=95680 225760 0 0 $X=95490 $Y=225520
X1635 VSS VDD ICV_23 $T=104420 29920 1 0 $X=104230 $Y=26960
X1636 VSS VDD ICV_23 $T=108100 198560 1 0 $X=107910 $Y=195600
X1637 VSS VDD ICV_23 $T=109480 149600 1 0 $X=109290 $Y=146640
X1638 VSS VDD ICV_23 $T=152260 13600 1 0 $X=152070 $Y=10640
X1639 VSS VDD ICV_23 $T=167900 144160 1 0 $X=167710 $Y=141200
X1640 VSS VDD ICV_23 $T=171580 165920 1 0 $X=171390 $Y=162960
X1641 VSS VDD ICV_23 $T=178480 46240 0 0 $X=178290 $Y=46000
X1642 VSS VDD ICV_23 $T=178480 149600 0 0 $X=178290 $Y=149360
X1643 VSS VDD ICV_23 $T=178940 29920 0 0 $X=178750 $Y=29680
X1644 VSS VDD ICV_23 $T=178940 106080 1 0 $X=178750 $Y=103120
X1645 VSS VDD ICV_23 $T=184460 111520 0 0 $X=184270 $Y=111280
X1646 VSS VDD ICV_23 $T=188600 160480 1 0 $X=188410 $Y=157520
X1647 VSS VDD ICV_23 $T=189060 40800 0 0 $X=188870 $Y=40560
X1648 VSS VDD ICV_23 $T=200100 138720 1 0 $X=199910 $Y=135760
X1649 VSS VDD ICV_23 $T=202400 149600 1 0 $X=202210 $Y=146640
X1650 VSS VDD ICV_23 $T=212060 68000 0 0 $X=211870 $Y=67760
X1651 VSS VDD ICV_23 $T=212060 220320 0 0 $X=211870 $Y=220080
X1652 VSS VDD ICV_24 $T=15640 209440 1 0 $X=15450 $Y=206480
X1653 VSS VDD ICV_24 $T=71760 46240 1 0 $X=71570 $Y=43280
X1654 VSS VDD ICV_24 $T=71760 100640 1 0 $X=71570 $Y=97680
X1655 VSS VDD ICV_24 $T=71760 111520 1 0 $X=71570 $Y=108560
X1656 VSS VDD ICV_24 $T=99820 160480 1 0 $X=99630 $Y=157520
X1657 VSS VDD ICV_24 $T=127880 138720 1 0 $X=127690 $Y=135760
X1658 VSS VDD ICV_24 $T=184000 24480 1 0 $X=183810 $Y=21520
X1659 VSS VDD ICV_24 $T=197800 198560 0 0 $X=197610 $Y=198320
X1660 VSS VDD ICV_24 $T=212060 46240 1 0 $X=211870 $Y=43280
X1661 VSS VDD ICV_24 $T=212060 182240 1 0 $X=211870 $Y=179280
X1662 VSS VDD 42 63 43 71 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=10120 73440 1 0 $X=9930 $Y=70480
X1663 VSS VDD 61 85 77 22 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=14260 40800 0 0 $X=14070 $Y=40560
X1664 VSS VDD 19 139 147 170 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=26680 24480 1 0 $X=26490 $Y=21520
X1665 VSS VDD 19 157 168 182 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=30360 46240 1 0 $X=30170 $Y=43280
X1666 VSS VDD 263 SCAN_IN<8> 271 292 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=50140 155040 1 0 $X=49950 $Y=152080
X1667 VSS VDD 58 343 470 457 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=91080 204000 1 0 $X=90890 $Y=201040
X1668 VSS VDD 58 535 642 621 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=120520 209440 1 0 $X=120330 $Y=206480
X1669 VSS VDD 706 708 671 663 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=133860 220320 0 0 $X=133670 $Y=220080
X1670 VSS VDD 679 SCAN_IN<8> 719 724 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=136160 13600 0 0 $X=135970 $Y=13360
X1671 VSS VDD 596 802 886 831 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=167900 73440 1 0 $X=167710 $Y=70480
X1672 VSS VDD 837 863 798 868 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=167900 209440 1 0 $X=167710 $Y=206480
X1673 VSS VDD 596 861 876 858 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=169280 122400 1 0 $X=169090 $Y=119440
X1674 VSS VDD 900 899 851 859 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=172960 133280 1 0 $X=172770 $Y=130320
X1675 VSS VDD 507 907 889 883 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=175260 204000 0 0 $X=175070 $Y=203760
X1676 VSS VDD 1005 984 727 1016 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=203780 165920 0 0 $X=203590 $Y=165680
X1677 VSS VDD 1012 SCAN_IN<1> 819 1023 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=206080 182240 1 0 $X=205890 $Y=179280
X1678 VSS VDD 1003 1025 1048 1032 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=212060 160480 0 0 $X=211870 $Y=160240
X1679 VSS VDD 19 53 72 VDD 21 VSS sky130_fd_sc_hd__nor3_4 $T=7820 24480 0 0 $X=7630 $Y=24240
X1680 VSS VDD 58 48 34 VDD 83 VSS sky130_fd_sc_hd__nor3_4 $T=8740 193120 0 0 $X=8550 $Y=192880
X1681 VSS VDD 19 22 54 VDD 23 VSS sky130_fd_sc_hd__nor3_4 $T=9660 46240 1 0 $X=9470 $Y=43280
X1682 VSS VDD 49 70 88 VDD 124 VSS sky130_fd_sc_hd__nor3_4 $T=16560 19040 0 0 $X=16370 $Y=18800
X1683 VSS VDD 19 167 163 VDD 178 VSS sky130_fd_sc_hd__nor3_4 $T=23920 29920 0 0 $X=23730 $Y=29680
X1684 VSS VDD 118 189 190 VDD 111 VSS sky130_fd_sc_hd__nor3_4 $T=33120 198560 1 0 $X=32930 $Y=195600
X1685 VSS VDD 92 208 197 VDD 202 VSS sky130_fd_sc_hd__nor3_4 $T=34040 214880 1 0 $X=33850 $Y=211920
X1686 VSS VDD 154 203 209 VDD 227 VSS sky130_fd_sc_hd__nor3_4 $T=35420 19040 0 0 $X=35230 $Y=18800
X1687 VSS VDD 231 240 245 VDD 208 VSS sky130_fd_sc_hd__nor3_4 $T=41400 204000 0 0 $X=41210 $Y=203760
X1688 VSS VDD 307 351 318 VDD 254 VSS sky130_fd_sc_hd__nor3_4 $T=59340 51680 1 0 $X=59150 $Y=48720
X1689 VSS VDD 339 189 190 VDD 313 VSS sky130_fd_sc_hd__nor3_4 $T=63020 193120 0 0 $X=62830 $Y=192880
X1690 VSS VDD 378 240 245 VDD 398 VSS sky130_fd_sc_hd__nor3_4 $T=70380 204000 0 0 $X=70190 $Y=203760
X1691 VSS VDD 460 240 245 VDD 462 VSS sky130_fd_sc_hd__nor3_4 $T=86480 209440 1 0 $X=86290 $Y=206480
X1692 VSS VDD 337 189 190 VDD 469 VSS sky130_fd_sc_hd__nor3_4 $T=89240 187680 1 0 $X=89050 $Y=184720
X1693 VSS VDD 507 240 245 VDD 541 VSS sky130_fd_sc_hd__nor3_4 $T=97060 209440 0 0 $X=96870 $Y=209200
X1694 VSS VDD 568 189 190 VDD 539 VSS sky130_fd_sc_hd__nor3_4 $T=108100 187680 0 0 $X=107910 $Y=187440
X1695 VSS VDD 596 606 572 VDD 527 VSS sky130_fd_sc_hd__nor3_4 $T=113160 68000 1 0 $X=112970 $Y=65040
X1696 VSS VDD 395 645 619 VDD 580 VSS sky130_fd_sc_hd__nor3_4 $T=116840 187680 1 0 $X=116650 $Y=184720
X1697 VSS VDD 620 189 190 VDD 626 VSS sky130_fd_sc_hd__nor3_4 $T=119140 193120 0 0 $X=118950 $Y=192880
X1698 VSS VDD 623 730 703 VDD 587 VSS sky130_fd_sc_hd__nor3_4 $T=133400 46240 1 0 $X=133210 $Y=43280
X1699 VSS VDD 551 754 740 VDD 735 VSS sky130_fd_sc_hd__nor3_4 $T=143060 46240 1 0 $X=142870 $Y=43280
X1700 VSS VDD 628 766 755 VDD 754 VSS sky130_fd_sc_hd__nor3_4 $T=146740 57120 1 0 $X=146550 $Y=54160
X1701 VSS VDD 756 766 755 VDD 803 VSS sky130_fd_sc_hd__nor3_4 $T=151340 68000 0 0 $X=151150 $Y=67760
X1702 VSS VDD 723 766 755 VDD 799 VSS sky130_fd_sc_hd__nor3_4 $T=151340 138720 0 0 $X=151150 $Y=138480
X1703 VSS VDD 757 766 755 VDD 813 VSS sky130_fd_sc_hd__nor3_4 $T=153640 133280 0 0 $X=153450 $Y=133040
X1704 VSS VDD 774 730 703 VDD 832 VSS sky130_fd_sc_hd__nor3_4 $T=159620 100640 0 0 $X=159430 $Y=100400
X1705 VSS VDD 830 730 703 VDD 805 VSS sky130_fd_sc_hd__nor3_4 $T=161460 46240 1 0 $X=161270 $Y=43280
X1706 VSS VDD 771 730 703 VDD 850 VSS sky130_fd_sc_hd__nor3_4 $T=161460 84320 1 0 $X=161270 $Y=81360
X1707 VSS VDD 776 730 703 VDD 856 VSS sky130_fd_sc_hd__nor3_4 $T=161460 106080 0 0 $X=161270 $Y=105840
X1708 VSS VDD 895 905 896 VDD 924 VSS sky130_fd_sc_hd__nor3_4 $T=185380 176800 0 0 $X=185190 $Y=176560
X1709 VSS VDD 980 990 968 VDD 952 VSS sky130_fd_sc_hd__nor3_4 $T=195500 220320 1 0 $X=195310 $Y=217360
X1710 VSS VDD 986 996 995 VDD 1009 VSS sky130_fd_sc_hd__nor3_4 $T=201480 89760 1 0 $X=201290 $Y=86800
X1711 VSS VDD 1004 1020 1028 VDD 818 VSS sky130_fd_sc_hd__nor3_4 $T=205620 19040 0 0 $X=205430 $Y=18800
X1712 VSS VDD 1007 1026 1023 VDD 1013 VSS sky130_fd_sc_hd__nor3_4 $T=206540 193120 1 0 $X=206350 $Y=190160
X1713 VSS VDD 1040 1045 1051 VDD 1028 VSS sky130_fd_sc_hd__nor3_4 $T=212060 24480 0 0 $X=211870 $Y=24240
X1714 VSS VDD 1041 1046 1050 VDD 1051 VSS sky130_fd_sc_hd__nor3_4 $T=212060 57120 0 0 $X=211870 $Y=56880
X1715 VSS VDD 1043 1042 1049 VDD 1050 VSS sky130_fd_sc_hd__nor3_4 $T=212060 149600 0 0 $X=211870 $Y=149360
X1716 VSS VDD 25 62 ICV_25 $T=10120 62560 1 0 $X=9930 $Y=59600
X1717 VSS VDD 153 80 ICV_25 $T=22080 51680 0 0 $X=21890 $Y=51440
X1718 VSS VDD 177 194 ICV_25 $T=36340 116960 1 0 $X=36150 $Y=114000
X1719 VSS VDD 386 412 ICV_25 $T=86480 24480 1 0 $X=86290 $Y=21520
X1720 VSS VDD 253 SCAN_IN<8> ICV_25 $T=90620 19040 1 0 $X=90430 $Y=16080
X1721 VSS VDD 476 377 ICV_25 $T=93840 155040 1 0 $X=93650 $Y=152080
X1722 VSS VDD 499 538 ICV_25 $T=105340 176800 1 0 $X=105150 $Y=173840
X1723 VSS VDD 512 618 ICV_25 $T=119140 165920 0 0 $X=118950 $Y=165680
X1724 VSS VDD 650 548 ICV_25 $T=122360 73440 0 0 $X=122170 $Y=73200
X1725 VSS VDD 733 SCAN_IN<12> ICV_25 $T=134780 133280 0 0 $X=134590 $Y=133040
X1726 VSS VDD 770 460 ICV_25 $T=143520 209440 1 0 $X=143330 $Y=206480
X1727 VSS VDD 772 753 ICV_25 $T=148580 127840 1 0 $X=148390 $Y=124880
X1728 VSS VDD 953 969 ICV_25 $T=196420 29920 1 0 $X=196230 $Y=26960
X1729 VSS VDD 998 723 ICV_25 $T=199180 155040 1 0 $X=198990 $Y=152080
X1730 VSS VDD 1019 SCAN_IN<4> ICV_25 $T=212060 100640 0 0 $X=211870 $Y=100400
X1731 VSS VDD 10 ICV_26 $T=33580 29920 1 0 $X=33390 $Y=26960
X1732 VSS VDD 10 ICV_26 $T=38180 51680 1 0 $X=37990 $Y=48720
X1733 VSS VDD 177 ICV_26 $T=44160 111520 0 0 $X=43970 $Y=111280
X1734 VSS VDD 331 ICV_26 $T=76360 144160 0 0 $X=76170 $Y=143920
X1735 VSS VDD 497 ICV_26 $T=94300 106080 1 0 $X=94110 $Y=103120
X1736 VSS VDD 326 ICV_26 $T=97520 100640 0 0 $X=97330 $Y=100400
X1737 VSS VDD 566 ICV_26 $T=106260 78880 0 0 $X=106070 $Y=78640
X1738 VSS VDD 579 ICV_26 $T=108100 111520 1 0 $X=107910 $Y=108560
X1739 VSS VDD 698 ICV_26 $T=132480 84320 0 0 $X=132290 $Y=84080
X1740 VSS VDD 703 ICV_26 $T=133400 40800 1 0 $X=133210 $Y=37840
X1741 VSS VDD 706 ICV_26 $T=133860 209440 1 0 $X=133670 $Y=206480
X1742 VSS VDD 768 ICV_26 $T=148580 95200 1 0 $X=148390 $Y=92240
X1743 VSS VDD 1002 ICV_26 $T=212060 89760 0 0 $X=211870 $Y=89520
X1744 VSS VDD 69 68 57 50 VDD 67 VSS sky130_fd_sc_hd__o22a_4 $T=9660 155040 0 0 $X=9470 $Y=154800
X1745 VSS VDD 105 130 173 SCAN_IN<10> VDD 82 VSS sky130_fd_sc_hd__o22a_4 $T=23920 149600 1 0 $X=23730 $Y=146640
X1746 VSS VDD 57 188 148 187 VDD 196 VSS sky130_fd_sc_hd__o22a_4 $T=30820 155040 1 0 $X=30630 $Y=152080
X1747 VSS VDD 87 118 127 231 VDD 213 VSS sky130_fd_sc_hd__o22a_4 $T=34960 193120 0 0 $X=34770 $Y=192880
X1748 VSS VDD 64 226 91 214 VDD 220 VSS sky130_fd_sc_hd__o22a_4 $T=36340 106080 1 0 $X=36150 $Y=103120
X1749 VSS VDD 263 252 258 253 VDD 68 VSS sky130_fd_sc_hd__o22a_4 $T=45080 155040 0 0 $X=44890 $Y=154800
X1750 VSS VDD 348 339 349 378 VDD 389 VSS sky130_fd_sc_hd__o22a_4 $T=69920 182240 0 0 $X=69730 $Y=182000
X1751 VSS VDD 425 407 348 418 VDD 252 VSS sky130_fd_sc_hd__o22a_4 $T=74520 155040 0 0 $X=74330 $Y=154800
X1752 VSS VDD 386 147 412 365 VDD 344 VSS sky130_fd_sc_hd__o22a_4 $T=77280 24480 1 0 $X=77090 $Y=21520
X1753 VSS VDD 389 385 395 424 VDD 426 VSS sky130_fd_sc_hd__o22a_4 $T=77280 187680 1 0 $X=77090 $Y=184720
X1754 VSS VDD 432 438 431 461 VDD 406 VSS sky130_fd_sc_hd__o22a_4 $T=82340 122400 0 0 $X=82150 $Y=122160
X1755 VSS VDD 449 230 413 188 VDD 436 VSS sky130_fd_sc_hd__o22a_4 $T=82800 133280 1 0 $X=82610 $Y=130320
X1756 VSS VDD 466 282 473 453 VDD 440 VSS sky130_fd_sc_hd__o22a_4 $T=87860 78880 1 0 $X=87670 $Y=75920
X1757 VSS VDD 466 415 473 454 VDD 427 VSS sky130_fd_sc_hd__o22a_4 $T=91080 78880 0 0 $X=90890 $Y=78640
X1758 VSS VDD 466 484 473 511 VDD 455 VSS sky130_fd_sc_hd__o22a_4 $T=95680 95200 0 0 $X=95490 $Y=94960
X1759 VSS VDD 533 516 522 50 VDD 508 VSS sky130_fd_sc_hd__o22a_4 $T=101660 19040 0 0 $X=101470 $Y=18800
X1760 VSS VDD 510 130 534 SCAN_IN<10> VDD 514 VSS sky130_fd_sc_hd__o22a_4 $T=101660 57120 0 0 $X=101470 $Y=56880
X1761 VSS VDD SCAN_IN<11> 471 SCAN_IN<12> 537 VDD 517 VSS sky130_fd_sc_hd__o22a_4 $T=105340 133280 0 0 $X=105150 $Y=133040
X1762 VSS VDD 466 579 346 592 VDD 296 VSS sky130_fd_sc_hd__o22a_4 $T=108100 116960 1 0 $X=107910 $Y=114000
X1763 VSS VDD 634 184 633 301 VDD 583 VSS sky130_fd_sc_hd__o22a_4 $T=117760 220320 1 0 $X=117570 $Y=217360
X1764 VSS VDD 522 628 604 632 VDD 649 VSS sky130_fd_sc_hd__o22a_4 $T=120980 51680 1 0 $X=120790 $Y=48720
X1765 VSS VDD 668 636 489 623 VDD 643 VSS sky130_fd_sc_hd__o22a_4 $T=121900 40800 1 0 $X=121710 $Y=37840
X1766 VSS VDD 672 449 666 413 VDD 648 VSS sky130_fd_sc_hd__o22a_4 $T=126500 106080 0 0 $X=126310 $Y=105840
X1767 VSS VDD 679 697 676 253 VDD 516 VSS sky130_fd_sc_hd__o22a_4 $T=133400 19040 1 0 $X=133210 $Y=16080
X1768 VSS VDD SCAN_IN<13> 680 693 673 VDD 472 VSS sky130_fd_sc_hd__o22a_4 $T=133400 144160 1 0 $X=133210 $Y=141200
X1769 VSS VDD 738 680 641 620 VDD 691 VSS sky130_fd_sc_hd__o22a_4 $T=139380 193120 1 0 $X=139190 $Y=190160
X1770 VSS VDD 753 743 737 732 VDD 746 VSS sky130_fd_sc_hd__o22a_4 $T=140760 122400 1 0 $X=140570 $Y=119440
X1771 VSS VDD 761 741 325 760 VDD 407 VSS sky130_fd_sc_hd__o22a_4 $T=144440 165920 1 0 $X=144250 $Y=162960
X1772 VSS VDD 748 773 676 628 VDD 668 VSS sky130_fd_sc_hd__o22a_4 $T=147200 35360 0 0 $X=147010 $Y=35120
X1773 VSS VDD 644 774 771 589 VDD 704 VSS sky130_fd_sc_hd__o22a_4 $T=147200 111520 1 0 $X=147010 $Y=108560
X1774 VSS VDD 757 758 776 693 VDD 753 VSS sky130_fd_sc_hd__o22a_4 $T=147200 127840 0 0 $X=147010 $Y=127600
X1775 VSS VDD 751 779 590 750 VDD 528 VSS sky130_fd_sc_hd__o22a_4 $T=147200 176800 0 0 $X=147010 $Y=176560
X1776 VSS VDD 778 763 690 680 VDD 751 VSS sky130_fd_sc_hd__o22a_4 $T=149500 187680 1 0 $X=149310 $Y=184720
X1777 VSS VDD 633 471 795 798 VDD 778 VSS sky130_fd_sc_hd__o22a_4 $T=155480 198560 0 0 $X=155290 $Y=198320
X1778 VSS VDD 759 677 819 745 VDD 785 VSS sky130_fd_sc_hd__o22a_4 $T=161460 144160 1 0 $X=161270 $Y=141200
X1779 VSS VDD 853 864 865 418 VDD 697 VSS sky130_fd_sc_hd__o22a_4 $T=167900 19040 1 0 $X=167710 $Y=16080
X1780 VSS VDD 883 857 624 873 VDD 841 VSS sky130_fd_sc_hd__o22a_4 $T=170200 198560 1 0 $X=170010 $Y=195600
X1781 VSS VDD 855 SCAN_IN<1> 634 917 VDD 863 VSS sky130_fd_sc_hd__o22a_4 $T=178940 220320 0 0 $X=178750 $Y=220080
X1782 VSS VDD 896 905 547 914 VDD 903 VSS sky130_fd_sc_hd__o22a_4 $T=179400 182240 0 0 $X=179210 $Y=182000
X1783 VSS VDD 769 723 759 940 VDD 943 VSS sky130_fd_sc_hd__o22a_4 $T=184920 144160 0 0 $X=184730 $Y=143920
X1784 VSS VDD 942 936 892 776 VDD 944 VSS sky130_fd_sc_hd__o22a_4 $T=185840 127840 0 0 $X=185650 $Y=127600
X1785 VSS VDD 943 939 851 757 VDD 942 VSS sky130_fd_sc_hd__o22a_4 $T=189520 138720 1 0 $X=189330 $Y=135760
X1786 VSS VDD 981 974 953 760 VDD 864 VSS sky130_fd_sc_hd__o22a_4 $T=194120 19040 1 0 $X=193930 $Y=16080
X1787 VSS VDD 982 971 927 988 VDD 964 VSS sky130_fd_sc_hd__o22a_4 $T=195500 116960 1 0 $X=195310 $Y=114000
X1788 VSS VDD 983 975 913 973 VDD 982 VSS sky130_fd_sc_hd__o22a_4 $T=195960 144160 1 0 $X=195770 $Y=141200
X1789 VSS VDD 819 661 928 727 VDD 983 VSS sky130_fd_sc_hd__o22a_4 $T=195960 149600 1 0 $X=195770 $Y=146640
X1790 VSS VDD 819 SCAN_IN<1> 915 917 VDD 984 VSS sky130_fd_sc_hd__o22a_4 $T=195960 182240 1 0 $X=195770 $Y=179280
X1791 VSS VDD 995 996 976 914 VDD 1002 VSS sky130_fd_sc_hd__o22a_4 $T=203320 95200 0 0 $X=203130 $Y=94960
X1792 VSS VDD 795 SCAN_IN<2> 671 1014 VDD 1011 VSS sky130_fd_sc_hd__o22a_4 $T=207920 214880 0 0 $X=207730 $Y=214640
X1793 VSS VDD 1023 1026 851 1014 VDD 1017 VSS sky130_fd_sc_hd__o22a_4 $T=209300 198560 0 0 $X=209110 $Y=198320
X1794 VSS VDD 1032 1052 988 1031 VDD 1049 VSS sky130_fd_sc_hd__o22a_4 $T=211600 155040 0 0 $X=211410 $Y=154800
X1795 VSS VDD 113 93 113 ICV_27 $T=19320 127840 0 0 $X=19130 $Y=127600
X1796 VSS VDD 91 152 91 ICV_27 $T=21620 106080 0 0 $X=21430 $Y=105840
X1797 VSS VDD 104 96 176 ICV_27 $T=23920 171360 0 0 $X=23730 $Y=171120
X1798 VSS VDD 138 280 138 ICV_27 $T=43240 220320 0 0 $X=43050 $Y=220080
X1799 VSS VDD 389 394 389 ICV_27 $T=69920 193120 0 0 $X=69730 $Y=192880
X1800 VSS VDD 365 390 365 ICV_27 $T=72680 13600 0 0 $X=72490 $Y=13360
X1801 VSS VDD 184 420 184 ICV_27 $T=73600 220320 0 0 $X=73410 $Y=220080
X1802 VSS VDD 493 502 493 ICV_27 $T=93380 40800 0 0 $X=93190 $Y=40560
X1803 VSS VDD 505 447 492 ICV_27 $T=94760 220320 0 0 $X=94570 $Y=220080
X1804 VSS VDD 525 554 525 ICV_27 $T=101200 13600 0 0 $X=101010 $Y=13360
X1805 VSS VDD 652 658 664 ICV_27 $T=122360 100640 1 0 $X=122170 $Y=97680
X1806 VSS VDD 635 651 635 ICV_27 $T=124200 171360 0 0 $X=124010 $Y=171120
X1807 VSS VDD 929 910 929 ICV_27 $T=181240 155040 0 0 $X=181050 $Y=154800
X1808 VSS VDD 926 921 926 ICV_27 $T=181700 84320 0 0 $X=181510 $Y=84080
X1809 VSS VDD SCAN_IN<4> 932 SCAN_IN<5> ICV_27 $T=188600 165920 0 0 $X=188410 $Y=165680
X1810 VSS VDD 945 976 945 ICV_27 $T=192280 100640 0 0 $X=192090 $Y=100400
X1811 VSS VDD SCAN_IN<1> 917 SCAN_IN<1> ICV_27 $T=195500 225760 0 0 $X=195310 $Y=225520
X1812 VSS VDD 987 1034 987 ICV_27 $T=208380 78880 0 0 $X=208190 $Y=78640
X1813 VSS VDD 1003 973 1003 ICV_27 $T=210220 144160 0 0 $X=210030 $Y=143920
X1814 VSS VDD SCAN_IN<2> 1014 SCAN_IN<2> ICV_27 $T=211140 209440 0 0 $X=210950 $Y=209200
X1815 VSS VDD 27 26 VDD 28 VSS sky130_fd_sc_hd__nand2_4 $T=7820 100640 1 0 $X=7630 $Y=97680
X1816 VSS VDD 29 37 VDD 36 VSS sky130_fd_sc_hd__nand2_4 $T=10120 89760 0 0 $X=9930 $Y=89520
X1817 VSS VDD 44 55 VDD 74 VSS sky130_fd_sc_hd__nand2_4 $T=10580 78880 0 0 $X=10390 $Y=78640
X1818 VSS VDD 257 247 VDD 278 VSS sky130_fd_sc_hd__nand2_4 $T=46460 122400 0 0 $X=46270 $Y=122160
X1819 VSS VDD 308 315 VDD 304 VSS sky130_fd_sc_hd__nand2_4 $T=54740 127840 0 0 $X=54550 $Y=127600
X1820 VSS VDD 363 347 VDD 358 VSS sky130_fd_sc_hd__nand2_4 $T=65320 138720 1 0 $X=65130 $Y=135760
X1821 VSS VDD 486 476 VDD 475 VSS sky130_fd_sc_hd__nand2_4 $T=92460 144160 1 0 $X=92270 $Y=141200
X1822 VSS VDD 561 568 VDD 486 VSS sky130_fd_sc_hd__nand2_4 $T=105340 149600 1 0 $X=105150 $Y=146640
X1823 VSS VDD 583 492 VDD 553 VSS sky130_fd_sc_hd__nand2_4 $T=108560 225760 1 0 $X=108370 $Y=222800
X1824 VSS VDD 290 634 VDD 582 VSS sky130_fd_sc_hd__nand2_4 $T=116380 225760 1 0 $X=116190 $Y=222800
X1825 VSS VDD 629 598 VDD 639 VSS sky130_fd_sc_hd__nand2_4 $T=120520 84320 0 0 $X=120330 $Y=84080
X1826 VSS VDD 670 637 VDD 688 VSS sky130_fd_sc_hd__nand2_4 $T=128800 62560 0 0 $X=128610 $Y=62320
X1827 VSS VDD 790 759 VDD 777 VSS sky130_fd_sc_hd__nand2_4 $T=152260 149600 1 0 $X=152070 $Y=146640
X1828 VSS VDD 785 791 VDD 794 VSS sky130_fd_sc_hd__nand2_4 $T=152260 155040 1 0 $X=152070 $Y=152080
X1829 VSS VDD 958 902 VDD 966 VSS sky130_fd_sc_hd__nand2_4 $T=194120 46240 0 0 $X=193930 $Y=46000
X1830 VSS VDD 1008 784 VDD 1000 VSS sky130_fd_sc_hd__nand2_4 $T=203320 57120 0 0 $X=203130 $Y=56880
X1831 VSS VDD 999 930 VDD 993 VSS sky130_fd_sc_hd__nand2_4 $T=203780 40800 1 0 $X=203590 $Y=37840
X1832 VSS VDD 1015 963 VDD 1006 VSS sky130_fd_sc_hd__nand2_4 $T=204240 68000 0 0 $X=204050 $Y=67760
X1833 VSS VDD 997 973 VDD 1039 VSS sky130_fd_sc_hd__nand2_4 $T=210220 138720 0 0 $X=210030 $Y=138480
X1834 VSS VDD 1035 988 VDD 1022 VSS sky130_fd_sc_hd__nand2_4 $T=211140 116960 0 0 $X=210950 $Y=116720
X1835 VSS VDD 57 188 173 187 VDD 219 VSS sky130_fd_sc_hd__a2bb2o_4 $T=34960 155040 0 0 $X=34770 $Y=154800
X1836 VSS VDD 59 222 102 215 VDD 248 VSS sky130_fd_sc_hd__a2bb2o_4 $T=36800 176800 0 0 $X=36610 $Y=176560
X1837 VSS VDD 266 37 266 37 VDD 341 VSS sky130_fd_sc_hd__a2bb2o_4 $T=55660 89760 1 0 $X=55470 $Y=86800
X1838 VSS VDD 26 285 55 276 VDD 342 VSS sky130_fd_sc_hd__a2bb2o_4 $T=57040 84320 1 0 $X=56850 $Y=81360
X1839 VSS VDD 330 119 26 285 VDD 360 VSS sky130_fd_sc_hd__a2bb2o_4 $T=58420 78880 1 0 $X=58230 $Y=75920
X1840 VSS VDD 325 337 258 324 VDD 329 VSS sky130_fd_sc_hd__a2bb2o_4 $T=59340 165920 1 0 $X=59150 $Y=162960
X1841 VSS VDD 334 326 345 326 VDD 154 VSS sky130_fd_sc_hd__a2bb2o_4 $T=63020 95200 0 0 $X=62830 $Y=94960
X1842 VSS VDD 371 374 396 399 VDD 411 VSS sky130_fd_sc_hd__a2bb2o_4 $T=68540 214880 0 0 $X=68350 $Y=214640
X1843 VSS VDD 128 383 373 168 VDD 369 VSS sky130_fd_sc_hd__a2bb2o_4 $T=69460 46240 0 0 $X=69270 $Y=46000
X1844 VSS VDD SCAN_IN<18> 315 422 388 VDD 439 VSS sky130_fd_sc_hd__a2bb2o_4 $T=74980 116960 0 0 $X=74790 $Y=116720
X1845 VSS VDD 407 429 407 429 VDD 364 VSS sky130_fd_sc_hd__a2bb2o_4 $T=78200 160480 0 0 $X=78010 $Y=160240
X1846 VSS VDD SCAN_IN<15> 512 589 377 VDD 575 VSS sky130_fd_sc_hd__a2bb2o_4 $T=105800 122400 1 0 $X=105610 $Y=119440
X1847 VSS VDD 590 512 481 337 VDD 640 VSS sky130_fd_sc_hd__a2bb2o_4 $T=115460 176800 1 0 $X=115270 $Y=173840
X1848 VSS VDD 522 623 519 637 VDD 636 VSS sky130_fd_sc_hd__a2bb2o_4 $T=120520 40800 0 0 $X=120330 $Y=40560
X1849 VSS VDD 654 595 647 576 VDD 683 VSS sky130_fd_sc_hd__a2bb2o_4 $T=122820 220320 0 0 $X=122630 $Y=220080
X1850 VSS VDD 522 628 534 632 VDD 695 VSS sky130_fd_sc_hd__a2bb2o_4 $T=125580 46240 0 0 $X=125390 $Y=46000
X1851 VSS VDD 590 750 752 507 VDD 779 VSS sky130_fd_sc_hd__a2bb2o_4 $T=145820 176800 1 0 $X=145630 $Y=173840
X1852 VSS VDD 749 SCAN_IN<18> 765 422 VDD 726 VSS sky130_fd_sc_hd__a2bb2o_4 $T=147200 84320 0 0 $X=147010 $Y=84080
X1853 VSS VDD 761 741 761 741 VDD 410 VSS sky130_fd_sc_hd__a2bb2o_4 $T=147200 165920 0 0 $X=147010 $Y=165680
X1854 VSS VDD 325 760 325 760 VDD 761 VSS sky130_fd_sc_hd__a2bb2o_4 $T=147660 160480 0 0 $X=147470 $Y=160240
X1855 VSS VDD 810 771 700 830 VDD 869 VSS sky130_fd_sc_hd__a2bb2o_4 $T=162840 35360 0 0 $X=162650 $Y=35120
X1856 VSS VDD 816 808 822 835 VDD 870 VSS sky130_fd_sc_hd__a2bb2o_4 $T=162840 127840 0 0 $X=162650 $Y=127600
X1857 VSS VDD 843 817 845 838 VDD 880 VSS sky130_fd_sc_hd__a2bb2o_4 $T=164680 68000 1 0 $X=164490 $Y=65040
X1858 VSS VDD 895 903 895 903 VDD 804 VSS sky130_fd_sc_hd__a2bb2o_4 $T=175260 176800 0 0 $X=175070 $Y=176560
X1859 VSS VDD 896 905 896 905 VDD 836 VSS sky130_fd_sc_hd__a2bb2o_4 $T=177100 187680 1 0 $X=176910 $Y=184720
X1860 VSS VDD 912 784 887 902 VDD 954 VSS sky130_fd_sc_hd__a2bb2o_4 $T=183080 51680 0 0 $X=182890 $Y=51440
X1861 VSS VDD 864 918 864 918 VDD 920 VSS sky130_fd_sc_hd__a2bb2o_4 $T=185380 13600 0 0 $X=185190 $Y=13360
X1862 VSS VDD 946 914 946 914 VDD 905 VSS sky130_fd_sc_hd__a2bb2o_4 $T=189520 182240 0 0 $X=189330 $Y=182000
X1863 VSS VDD 892 776 928 973 VDD 936 VSS sky130_fd_sc_hd__a2bb2o_4 $T=190440 133280 1 0 $X=190250 $Y=130320
X1864 VSS VDD 927 972 967 757 VDD 971 VSS sky130_fd_sc_hd__a2bb2o_4 $T=195040 122400 1 0 $X=194850 $Y=119440
X1865 VSS VDD 953 935 953 760 VDD 981 VSS sky130_fd_sc_hd__a2bb2o_4 $T=195500 24480 1 0 $X=195310 $Y=21520
X1866 VSS VDD 980 992 980 992 VDD 834 VSS sky130_fd_sc_hd__a2bb2o_4 $T=199640 209440 1 0 $X=199450 $Y=206480
X1867 VSS VDD 986 1002 986 1002 VDD 1037 VSS sky130_fd_sc_hd__a2bb2o_4 $T=203780 89760 0 0 $X=203590 $Y=89520
X1868 VSS VDD 976 1019 976 914 VDD 996 VSS sky130_fd_sc_hd__a2bb2o_4 $T=205160 100640 1 0 $X=204970 $Y=97680
X1869 VSS VDD 1023 1026 1023 1026 VDD 1048 VSS sky130_fd_sc_hd__a2bb2o_4 $T=210680 182240 0 0 $X=210490 $Y=182000
X1870 VSS VDD 1033 1014 1033 1014 VDD 1026 VSS sky130_fd_sc_hd__a2bb2o_4 $T=210680 204000 0 0 $X=210490 $Y=203760
X1871 VSS VDD 134 ICV_28 $T=20240 40800 1 0 $X=20050 $Y=37840
X1872 VSS VDD 138 ICV_28 $T=20240 220320 1 0 $X=20050 $Y=217360
X1873 VSS VDD 182 ICV_28 $T=27600 51680 1 0 $X=27410 $Y=48720
X1874 VSS VDD 211 ICV_28 $T=33120 84320 1 0 $X=32930 $Y=81360
X1875 VSS VDD 43 ICV_28 $T=34040 62560 0 0 $X=33850 $Y=62320
X1876 VSS VDD 242 ICV_28 $T=39560 95200 0 0 $X=39370 $Y=94960
X1877 VSS VDD 249 ICV_28 $T=42320 187680 0 0 $X=42130 $Y=187440
X1878 VSS VDD 294 ICV_28 $T=48300 35360 1 0 $X=48110 $Y=32400
X1879 VSS VDD 345 ICV_28 $T=59800 95200 1 0 $X=59610 $Y=92240
X1880 VSS VDD 326 ICV_28 $T=59800 100640 1 0 $X=59610 $Y=97680
X1881 VSS VDD CLK_OUT ICV_28 $T=67160 100640 0 0 $X=66970 $Y=100400
X1882 VSS VDD 400 ICV_28 $T=69920 149600 0 0 $X=69730 $Y=149360
X1883 VSS VDD 348 ICV_28 $T=70380 155040 0 0 $X=70190 $Y=154800
X1884 VSS VDD 632 ICV_28 $T=116840 51680 1 0 $X=116650 $Y=48720
X1885 VSS VDD 548 ICV_28 $T=118220 73440 0 0 $X=118030 $Y=73200
X1886 VSS VDD 637 ICV_28 $T=124660 62560 0 0 $X=124470 $Y=62320
X1887 VSS VDD 676 ICV_28 $T=126040 29920 0 0 $X=125850 $Y=29680
X1888 VSS VDD SCAN_IN<11> ICV_28 $T=126040 127840 0 0 $X=125850 $Y=127600
X1889 VSS VDD 653 ICV_28 $T=130640 182240 0 0 $X=130450 $Y=182000
X1890 VSS VDD 715 ICV_28 $T=132480 182240 1 0 $X=132290 $Y=179280
X1891 VSS VDD 578 ICV_28 $T=134780 57120 0 0 $X=134590 $Y=56880
X1892 VSS VDD 766 ICV_28 $T=144440 51680 1 0 $X=144250 $Y=48720
X1893 VSS VDD 782 ICV_28 $T=149040 46240 1 0 $X=148850 $Y=43280
X1894 VSS VDD 16 ICV_28 $T=149960 214880 0 0 $X=149770 $Y=214640
X1895 VSS VDD 592 ICV_28 $T=153640 116960 0 0 $X=153450 $Y=116720
X1896 VSS VDD 558 ICV_28 $T=161920 198560 0 0 $X=161730 $Y=198320
X1897 VSS VDD 966 ICV_28 $T=190900 51680 1 0 $X=190710 $Y=48720
X1898 VSS VDD 929 ICV_28 $T=192740 155040 0 0 $X=192550 $Y=154800
X1899 VSS VDD 701 ICV_28 $T=199640 40800 1 0 $X=199450 $Y=37840
X1900 VSS VDD 1008 ICV_28 $T=199640 57120 1 0 $X=199450 $Y=54160
X1901 VSS VDD 1013 ICV_28 $T=201940 187680 1 0 $X=201750 $Y=184720
X1902 VSS VDD 1034 ICV_28 $T=207000 73440 1 0 $X=206810 $Y=70480
X1903 VSS VDD SCAN_IN<17> ICV_28 $T=209760 95200 0 0 $X=209570 $Y=94960
X1904 VSS VDD 1048 ICV_28 $T=209760 165920 0 0 $X=209570 $Y=165680
X1905 VSS VDD 70 88 ICV_29 $T=11040 19040 0 0 $X=10850 $Y=18800
X1906 VSS VDD 117 128 ICV_29 $T=18400 29920 0 0 $X=18210 $Y=29680
X1907 VSS VDD 133 147 ICV_29 $T=22540 19040 1 0 $X=22350 $Y=16080
X1908 VSS VDD 33 149 ICV_29 $T=23000 176800 0 0 $X=22810 $Y=176560
X1909 VSS VDD 188 200 ICV_29 $T=29440 160480 1 0 $X=29250 $Y=157520
X1910 VSS VDD 212 20 ICV_29 $T=34040 116960 0 0 $X=33850 $Y=116720
X1911 VSS VDD 244 256 ICV_29 $T=40480 165920 0 0 $X=40290 $Y=165680
X1912 VSS VDD 297 310 ICV_29 $T=49220 220320 0 0 $X=49030 $Y=220080
X1913 VSS VDD 16 20 ICV_29 $T=50600 187680 0 0 $X=50410 $Y=187440
X1914 VSS VDD 313 320 ICV_29 $T=52440 198560 1 0 $X=52250 $Y=195600
X1915 VSS VDD 328 335 ICV_29 $T=56120 155040 1 0 $X=55930 $Y=152080
X1916 VSS VDD 430 430 ICV_29 $T=77280 24480 0 0 $X=77090 $Y=24240
X1917 VSS VDD 363 295 ICV_29 $T=84180 133280 0 0 $X=83990 $Y=133040
X1918 VSS VDD 474 299 ICV_29 $T=87860 116960 1 0 $X=87670 $Y=114000
X1919 VSS VDD 719 679 ICV_29 $T=134320 13600 1 0 $X=134130 $Y=10640
X1920 VSS VDD 721 733 ICV_29 $T=134320 127840 0 0 $X=134130 $Y=127600
X1921 VSS VDD 721 733 ICV_29 $T=137540 122400 0 0 $X=137350 $Y=122160
X1922 VSS VDD 775 780 ICV_29 $T=146740 29920 1 0 $X=146550 $Y=26960
X1923 VSS VDD 860 672 ICV_29 $T=165600 100640 0 0 $X=165410 $Y=100400
X1924 VSS VDD 865 756 ICV_29 $T=174340 29920 0 0 $X=174150 $Y=29680
X1925 VSS VDD SCAN_IN<3> SCAN_IN<2> ICV_29 $T=181700 209440 0 0 $X=181510 $Y=209200
X1926 VSS VDD 661 727 ICV_29 $T=202400 138720 0 0 $X=202210 $Y=138480
X1927 VSS VDD 1014 671 ICV_29 $T=202400 209440 0 0 $X=202210 $Y=209200
X1928 VSS VDD 795 SCAN_IN<2> ICV_29 $T=202400 214880 0 0 $X=202210 $Y=214640
X1929 VSS VDD 158 997 ICV_29 $T=207000 133280 1 0 $X=206810 $Y=130320
X1930 VSS VDD 1031 1052 ICV_29 $T=209760 160480 1 0 $X=209570 $Y=157520
X1931 VSS VDD 35 61 ICV_30 $T=6900 19040 0 0 $X=6710 $Y=18800
X1932 VSS VDD 40 65 ICV_30 $T=6900 187680 0 0 $X=6710 $Y=187440
X1933 VSS VDD 71 42 ICV_30 $T=11040 68000 1 0 $X=10850 $Y=65040
X1934 VSS VDD 79 127 ICV_30 $T=18400 214880 0 0 $X=18210 $Y=214640
X1935 VSS VDD 176 59 ICV_30 $T=31280 176800 1 0 $X=31090 $Y=173840
X1936 VSS VDD 20 202 ICV_30 $T=31280 220320 1 0 $X=31090 $Y=217360
X1937 VSS VDD 214 91 ICV_30 $T=34960 100640 1 0 $X=34770 $Y=97680
X1938 VSS VDD 57 187 ICV_30 $T=36340 165920 0 0 $X=36150 $Y=165680
X1939 VSS VDD 247 257 ICV_30 $T=41400 122400 0 0 $X=41210 $Y=122160
X1940 VSS VDD 356 348 ICV_30 $T=62100 155040 0 0 $X=61910 $Y=154800
X1941 VSS VDD 381 384 ICV_30 $T=67620 111520 1 0 $X=67430 $Y=108560
X1942 VSS VDD 330 289 ICV_30 $T=74980 51680 0 0 $X=74790 $Y=51440
X1943 VSS VDD 20 427 ICV_30 $T=75900 68000 0 0 $X=75710 $Y=67760
X1944 VSS VDD 416 20 ICV_30 $T=81420 89760 0 0 $X=81230 $Y=89520
X1945 VSS VDD 447 401 ICV_30 $T=82800 214880 0 0 $X=82610 $Y=214640
X1946 VSS VDD 16 480 ICV_30 $T=88780 176800 1 0 $X=88590 $Y=173840
X1947 VSS VDD 471 SCAN_IN<11> ICV_30 $T=100280 133280 0 0 $X=100090 $Y=133040
X1948 VSS VDD 478 575 ICV_30 $T=104420 122400 0 0 $X=104230 $Y=122160
X1949 VSS VDD 602 58 ICV_30 $T=110860 204000 0 0 $X=110670 $Y=203760
X1950 VSS VDD 610 109 ICV_30 $T=112700 155040 0 0 $X=112510 $Y=154800
X1951 VSS VDD 607 643 ICV_30 $T=117760 57120 1 0 $X=117570 $Y=54160
X1952 VSS VDD 625 620 ICV_30 $T=121440 155040 1 0 $X=121250 $Y=152080
X1953 VSS VDD 550 535 ICV_30 $T=121440 204000 1 0 $X=121250 $Y=201040
X1954 VSS VDD 665 620 ICV_30 $T=122820 187680 1 0 $X=122630 $Y=184720
X1955 VSS VDD 678 558 ICV_30 $T=126960 155040 0 0 $X=126770 $Y=154800
X1956 VSS VDD 537 690 ICV_30 $T=126960 187680 1 0 $X=126770 $Y=184720
X1957 VSS VDD 17 20 ICV_30 $T=134320 24480 0 0 $X=134130 $Y=24240
X1958 VSS VDD 747 460 ICV_30 $T=140300 204000 0 0 $X=140110 $Y=203760
X1959 VSS VDD 763 680 ICV_30 $T=144440 187680 1 0 $X=144250 $Y=184720
X1960 VSS VDD 731 755 ICV_30 $T=148580 73440 1 0 $X=148390 $Y=70480
X1961 VSS VDD 633 471 ICV_30 $T=154100 198560 1 0 $X=153910 $Y=195600
X1962 VSS VDD 513 815 ICV_30 $T=155940 46240 0 0 $X=155750 $Y=46000
X1963 VSS VDD 759 819 ICV_30 $T=157320 138720 0 0 $X=157130 $Y=138480
X1964 VSS VDD 17 20 ICV_30 $T=159160 24480 0 0 $X=158970 $Y=24240
X1965 VSS VDD 783 813 ICV_30 $T=159160 122400 0 0 $X=158970 $Y=122160
X1966 VSS VDD 863 837 ICV_30 $T=166520 204000 1 0 $X=166330 $Y=201040
X1967 VSS VDD 905 914 ICV_30 $T=174340 182240 0 0 $X=174150 $Y=182000
X1968 VSS VDD 889 907 ICV_30 $T=174340 198560 0 0 $X=174150 $Y=198320
X1969 VSS VDD 917 SCAN_IN<6> ICV_30 $T=177100 220320 1 0 $X=176910 $Y=217360
X1970 VSS VDD 922 888 ICV_30 $T=178480 95200 0 0 $X=178290 $Y=94960
X1971 VSS VDD 923 919 ICV_30 $T=178940 111520 1 0 $X=178750 $Y=108560
X1972 VSS VDD 910 723 ICV_30 $T=179860 144160 0 0 $X=179670 $Y=143920
X1973 VSS VDD 774 848 ICV_30 $T=187220 100640 0 0 $X=187030 $Y=100400
X1974 VSS VDD 953 760 ICV_30 $T=192740 13600 0 0 $X=192550 $Y=13360
X1975 VSS VDD 967 965 ICV_30 $T=195040 187680 0 0 $X=194850 $Y=187440
X1976 VSS VDD 991 998 ICV_30 $T=196420 160480 0 0 $X=196230 $Y=160240
X1977 VSS VDD 999 994 ICV_30 $T=199180 51680 1 0 $X=198990 $Y=48720
X1978 VSS VDD 985 20 ICV_30 $T=202400 111520 0 0 $X=202210 $Y=111280
X1979 VSS VDD 1026 1023 ICV_30 $T=205160 187680 1 0 $X=204970 $Y=184720
X1980 VSS VDD 1026 1023 ICV_30 $T=209300 187680 1 0 $X=209110 $Y=184720
X1981 VSS VDD 1033 851 ICV_30 $T=209300 204000 1 0 $X=209110 $Y=201040
X1982 VSS VDD 10 ICV_31 $T=21160 84320 1 0 $X=20970 $Y=81360
X1983 VSS VDD 209 ICV_31 $T=35420 24480 0 0 $X=35230 $Y=24240
X1984 VSS VDD 223 ICV_31 $T=49680 57120 0 0 $X=49490 $Y=56880
X1985 VSS VDD 284 ICV_31 $T=49680 62560 1 0 $X=49490 $Y=59600
X1986 VSS VDD 352 ICV_31 $T=63020 116960 1 0 $X=62830 $Y=114000
X1987 VSS VDD 20 ICV_31 $T=90160 182240 1 0 $X=89970 $Y=179280
X1988 VSS VDD SCAN_IN<8> ICV_31 $T=92460 13600 1 0 $X=92270 $Y=10640
X1989 VSS VDD 377 ICV_31 $T=94300 160480 0 0 $X=94110 $Y=160240
X1990 VSS VDD 672 ICV_31 $T=133400 89760 1 0 $X=133210 $Y=86800
X1991 VSS VDD 871 ICV_31 $T=174800 155040 1 0 $X=174610 $Y=152080
X1992 VSS VDD 834 ICV_31 $T=175720 187680 0 0 $X=175530 $Y=187440
X1993 VSS VDD 896 ICV_31 $T=189520 176800 1 0 $X=189330 $Y=173840
X1994 VSS VDD 1007 ICV_31 $T=209300 187680 0 0 $X=209110 $Y=187440
X1995 VSS VDD 33 79 VDD 65 VSS sky130_fd_sc_hd__and2_4 $T=12420 209440 1 0 $X=12230 $Y=206480
X1996 VSS VDD 49 88 VDD 72 VSS sky130_fd_sc_hd__and2_4 $T=17020 24480 0 0 $X=16830 $Y=24240
X1997 VSS VDD 59 106 VDD 40 VSS sky130_fd_sc_hd__and2_4 $T=18400 193120 0 0 $X=18210 $Y=192880
X1998 VSS VDD 114 93 VDD 137 VSS sky130_fd_sc_hd__and2_4 $T=20240 133280 0 0 $X=20050 $Y=133040
X1999 VSS VDD 87 106 VDD 97 VSS sky130_fd_sc_hd__and2_4 $T=20700 198560 0 0 $X=20510 $Y=198320
X2000 VSS VDD 87 115 VDD 141 VSS sky130_fd_sc_hd__and2_4 $T=21160 209440 1 0 $X=20970 $Y=206480
X2001 VSS VDD 128 88 VDD 163 VSS sky130_fd_sc_hd__and2_4 $T=24380 40800 1 0 $X=24190 $Y=37840
X2002 VSS VDD 153 193 VDD 204 VSS sky130_fd_sc_hd__and2_4 $T=34960 57120 0 0 $X=34770 $Y=56880
X2003 VSS VDD 57 187 VDD 237 VSS sky130_fd_sc_hd__and2_4 $T=37720 171360 1 0 $X=37530 $Y=168400
X2004 VSS VDD 127 225 VDD 197 VSS sky130_fd_sc_hd__and2_4 $T=37720 209440 0 0 $X=37530 $Y=209200
X2005 VSS VDD 177 226 VDD 217 VSS sky130_fd_sc_hd__and2_4 $T=40020 111520 0 0 $X=39830 $Y=111280
X2006 VSS VDD 258 253 VDD 263 VSS sky130_fd_sc_hd__and2_4 $T=48760 149600 0 0 $X=48570 $Y=149360
X2007 VSS VDD 127 231 VDD 300 VSS sky130_fd_sc_hd__and2_4 $T=49220 198560 1 0 $X=49030 $Y=195600
X2008 VSS VDD 310 297 VDD 305 VSS sky130_fd_sc_hd__and2_4 $T=54740 220320 0 0 $X=54550 $Y=220080
X2009 VSS VDD 84 312 VDD 287 VSS sky130_fd_sc_hd__and2_4 $T=57040 29920 1 0 $X=56850 $Y=26960
X2010 VSS VDD 310 106 VDD 320 VSS sky130_fd_sc_hd__and2_4 $T=57500 209440 1 0 $X=57310 $Y=206480
X2011 VSS VDD 348 356 VDD 336 VSS sky130_fd_sc_hd__and2_4 $T=67160 155040 0 0 $X=66970 $Y=154800
X2012 VSS VDD 310 339 VDD 385 VSS sky130_fd_sc_hd__and2_4 $T=67160 193120 1 0 $X=66970 $Y=190160
X2013 VSS VDD 372 350 VDD 318 VSS sky130_fd_sc_hd__and2_4 $T=68540 46240 1 0 $X=68350 $Y=43280
X2014 VSS VDD 275 43 VDD 387 VSS sky130_fd_sc_hd__and2_4 $T=69000 73440 1 0 $X=68810 $Y=70480
X2015 VSS VDD 349 290 VDD 396 VSS sky130_fd_sc_hd__and2_4 $T=69000 220320 1 0 $X=68810 $Y=217360
X2016 VSS VDD 390 376 VDD 382 VSS sky130_fd_sc_hd__and2_4 $T=72220 19040 0 0 $X=72030 $Y=18800
X2017 VSS VDD 345 7 VDD 367 VSS sky130_fd_sc_hd__and2_4 $T=77280 100640 1 0 $X=77090 $Y=97680
X2018 VSS VDD 413 231 VDD 428 VSS sky130_fd_sc_hd__and2_4 $T=78200 138720 1 0 $X=78010 $Y=135760
X2019 VSS VDD 420 437 VDD 442 VSS sky130_fd_sc_hd__and2_4 $T=80040 220320 1 0 $X=79850 $Y=217360
X2020 VSS VDD 464 442 VDD 477 VSS sky130_fd_sc_hd__and2_4 $T=87400 225760 1 0 $X=87210 $Y=222800
X2021 VSS VDD 464 290 VDD 483 VSS sky130_fd_sc_hd__and2_4 $T=91080 214880 0 0 $X=90890 $Y=214640
X2022 VSS VDD 481 106 VDD 446 VSS sky130_fd_sc_hd__and2_4 $T=92920 193120 0 0 $X=92730 $Y=192880
X2023 VSS VDD 554 50 VDD 533 VSS sky130_fd_sc_hd__and2_4 $T=105340 19040 1 0 $X=105150 $Y=16080
X2024 VSS VDD SCAN_IN<12> 537 VDD 494 VSS sky130_fd_sc_hd__and2_4 $T=108560 138720 1 0 $X=108370 $Y=135760
X2025 VSS VDD 489 574 VDD 593 VSS sky130_fd_sc_hd__and2_4 $T=110860 40800 0 0 $X=110670 $Y=40560
X2026 VSS VDD 529 591 VDD 606 VSS sky130_fd_sc_hd__and2_4 $T=110860 62560 0 0 $X=110670 $Y=62320
X2027 VSS VDD 507 549 VDD 625 VSS sky130_fd_sc_hd__and2_4 $T=118220 155040 1 0 $X=118030 $Y=152080
X2028 VSS VDD 641 290 VDD 627 VSS sky130_fd_sc_hd__and2_4 $T=122820 209440 0 0 $X=122630 $Y=209200
X2029 VSS VDD 489 657 VDD 609 VSS sky130_fd_sc_hd__and2_4 $T=125120 35360 1 0 $X=124930 $Y=32400
X2030 VSS VDD 700 253 VDD 679 VSS sky130_fd_sc_hd__and2_4 $T=133400 19040 0 0 $X=133210 $Y=18800
X2031 VSS VDD 633 537 VDD 665 VSS sky130_fd_sc_hd__and2_4 $T=133400 193120 1 0 $X=133210 $Y=190160
X2032 VSS VDD 676 744 VDD 740 VSS sky130_fd_sc_hd__and2_4 $T=147200 40800 0 0 $X=147010 $Y=40560
X2033 VSS VDD 776 693 VDD 743 VSS sky130_fd_sc_hd__and2_4 $T=150880 122400 1 0 $X=150690 $Y=119440
X2034 VSS VDD 788 574 VDD 797 VSS sky130_fd_sc_hd__and2_4 $T=153180 46240 1 0 $X=152990 $Y=43280
X2035 VSS VDD 738 798 VDD 763 VSS sky130_fd_sc_hd__and2_4 $T=161460 193120 1 0 $X=161270 $Y=190160
X2036 VSS VDD 851 790 VDD 822 VSS sky130_fd_sc_hd__and2_4 $T=166060 133280 1 0 $X=165870 $Y=130320
X2037 VSS VDD 810 790 VDD 845 VSS sky130_fd_sc_hd__and2_4 $T=168820 62560 1 0 $X=168630 $Y=59600
X2038 VSS VDD 892 790 VDD 849 VSS sky130_fd_sc_hd__and2_4 $T=175260 116960 0 0 $X=175070 $Y=116720
X2039 VSS VDD 769 894 VDD 852 VSS sky130_fd_sc_hd__and2_4 $T=175260 149600 0 0 $X=175070 $Y=149360
X2040 VSS VDD 759 721 VDD 939 VSS sky130_fd_sc_hd__and2_4 $T=185380 138720 0 0 $X=185190 $Y=138480
X2041 VSS VDD 929 SCAN_IN<0> VDD 978 VSS sky130_fd_sc_hd__and2_4 $T=192740 165920 1 0 $X=192550 $Y=162960
X2042 VSS VDD 928 727 VDD 975 VSS sky130_fd_sc_hd__and2_4 $T=195040 144160 0 0 $X=194850 $Y=143920
X2043 VSS VDD 904 920 VDD 1004 VSS sky130_fd_sc_hd__and2_4 $T=198260 13600 1 0 $X=198070 $Y=10640
X2044 VSS VDD 978 984 VDD 1012 VSS sky130_fd_sc_hd__and2_4 $T=201480 176800 1 0 $X=201290 $Y=173840
X2045 VSS VDD 1024 1036 VDD 1040 VSS sky130_fd_sc_hd__and2_4 $T=209300 24480 1 0 $X=209110 $Y=21520
X2046 VSS VDD 1034 1038 VDD 1042 VSS sky130_fd_sc_hd__and2_4 $T=209300 78880 1 0 $X=209110 $Y=75920
X2047 VSS VDD 988 1031 VDD 1043 VSS sky130_fd_sc_hd__and2_4 $T=209300 155040 1 0 $X=209110 $Y=152080
X2048 VSS VDD 44 55 VDD 63 VSS sky130_fd_sc_hd__or2_4 $T=11500 84320 1 0 $X=11310 $Y=81360
X2049 VSS VDD 73 80 VDD 77 VSS sky130_fd_sc_hd__or2_4 $T=12880 51680 1 0 $X=12690 $Y=48720
X2050 VSS VDD 25 91 VDD 66 VSS sky130_fd_sc_hd__or2_4 $T=15180 100640 0 0 $X=14990 $Y=100400
X2051 VSS VDD 101 110 VDD 20 VSS sky130_fd_sc_hd__or2_4 $T=21160 225760 1 0 $X=20970 $Y=222800
X2052 VSS VDD 149 33 VDD 143 VSS sky130_fd_sc_hd__or2_4 $T=24840 182240 1 0 $X=24650 $Y=179280
X2053 VSS VDD 133 61 VDD 139 VSS sky130_fd_sc_hd__or2_4 $T=25300 24480 0 0 $X=25110 $Y=24240
X2054 VSS VDD 181 164 VDD 198 VSS sky130_fd_sc_hd__or2_4 $T=29900 73440 1 0 $X=29710 $Y=70480
X2055 VSS VDD 175 136 VDD 160 VSS sky130_fd_sc_hd__or2_4 $T=31740 127840 1 0 $X=31550 $Y=124880
X2056 VSS VDD 117 128 VDD 133 VSS sky130_fd_sc_hd__or2_4 $T=34960 35360 0 0 $X=34770 $Y=35120
X2057 VSS VDD 136 SCAN_IN<20> VDD 228 VSS sky130_fd_sc_hd__or2_4 $T=36340 138720 0 0 $X=36150 $Y=138480
X2058 VSS VDD 206 161 VDD 225 VSS sky130_fd_sc_hd__or2_4 $T=36340 204000 1 0 $X=36150 $Y=201040
X2059 VSS VDD 238 279 VDD 259 VSS sky130_fd_sc_hd__or2_4 $T=48760 19040 0 0 $X=48570 $Y=18800
X2060 VSS VDD 256 188 VDD 268 VSS sky130_fd_sc_hd__or2_4 $T=49220 165920 1 0 $X=49030 $Y=162960
X2061 VSS VDD 286 271 VDD 149 VSS sky130_fd_sc_hd__or2_4 $T=50140 182240 0 0 $X=49950 $Y=182000
X2062 VSS VDD 242 266 VDD 267 VSS sky130_fd_sc_hd__or2_4 $T=51060 95200 1 0 $X=50870 $Y=92240
X2063 VSS VDD 267 276 VDD 284 VSS sky130_fd_sc_hd__or2_4 $T=51520 78880 0 0 $X=51330 $Y=78640
X2064 VSS VDD 359 166 VDD 371 VSS sky130_fd_sc_hd__or2_4 $T=64400 225760 1 0 $X=64210 $Y=222800
X2065 VSS VDD 363 347 VDD 308 VSS sky130_fd_sc_hd__or2_4 $T=65320 138720 0 0 $X=65130 $Y=138480
X2066 VSS VDD 379 373 VDD 391 VSS sky130_fd_sc_hd__or2_4 $T=80500 46240 0 0 $X=80310 $Y=46000
X2067 VSS VDD 391 383 VDD 430 VSS sky130_fd_sc_hd__or2_4 $T=82340 35360 1 0 $X=82150 $Y=32400
X2068 VSS VDD 430 412 VDD 238 VSS sky130_fd_sc_hd__or2_4 $T=82800 24480 0 0 $X=82610 $Y=24240
X2069 VSS VDD 486 476 VDD 363 VSS sky130_fd_sc_hd__or2_4 $T=92460 144160 0 0 $X=92270 $Y=143920
X2070 VSS VDD 442 464 VDD 505 VSS sky130_fd_sc_hd__or2_4 $T=92460 225760 0 0 $X=92270 $Y=225520
X2071 VSS VDD 538 506 VDD 433 VSS sky130_fd_sc_hd__or2_4 $T=105340 182240 1 0 $X=105150 $Y=179280
X2072 VSS VDD 629 598 VDD 562 VSS sky130_fd_sc_hd__or2_4 $T=119140 84320 1 0 $X=118950 $Y=81360
X2073 VSS VDD 476 SCAN_IN<16> VDD 630 VSS sky130_fd_sc_hd__or2_4 $T=119140 138720 0 0 $X=118950 $Y=138480
X2074 VSS VDD SCAN_IN<19> 637 VDD 656 VSS sky130_fd_sc_hd__or2_4 $T=120520 73440 1 0 $X=120330 $Y=70480
X2075 VSS VDD 624 SCAN_IN<14> VDD 531 VSS sky130_fd_sc_hd__or2_4 $T=123280 133280 1 0 $X=123090 $Y=130320
X2076 VSS VDD 670 637 VDD 629 VSS sky130_fd_sc_hd__or2_4 $T=127880 68000 0 0 $X=127690 $Y=67760
X2077 VSS VDD 674 676 VDD 657 VSS sky130_fd_sc_hd__or2_4 $T=131100 24480 0 0 $X=130910 $Y=24240
X2078 VSS VDD 706 690 VDD 642 VSS sky130_fd_sc_hd__or2_4 $T=133860 214880 1 0 $X=133670 $Y=211920
X2079 VSS VDD 713 690 VDD 550 VSS sky130_fd_sc_hd__or2_4 $T=137080 198560 1 0 $X=136890 $Y=195600
X2080 VSS VDD 437 734 VDD 708 VSS sky130_fd_sc_hd__or2_4 $T=137540 220320 1 0 $X=137350 $Y=217360
X2081 VSS VDD 464 634 VDD 734 VSS sky130_fd_sc_hd__or2_4 $T=143520 225760 1 0 $X=143330 $Y=222800
X2082 VSS VDD 747 633 VDD 728 VSS sky130_fd_sc_hd__or2_4 $T=147200 204000 0 0 $X=147010 $Y=203760
X2083 VSS VDD 770 747 VDD 786 VSS sky130_fd_sc_hd__or2_4 $T=153180 209440 1 0 $X=152990 $Y=206480
X2084 VSS VDD 796 788 VDD 789 VSS sky130_fd_sc_hd__or2_4 $T=155940 24480 0 0 $X=155750 $Y=24240
X2085 VSS VDD 799 783 VDD 814 VSS sky130_fd_sc_hd__or2_4 $T=156400 144160 0 0 $X=156210 $Y=143920
X2086 VSS VDD 803 783 VDD 838 VSS sky130_fd_sc_hd__or2_4 $T=161460 73440 1 0 $X=161270 $Y=70480
X2087 VSS VDD 813 783 VDD 835 VSS sky130_fd_sc_hd__or2_4 $T=161460 127840 1 0 $X=161270 $Y=124880
X2088 VSS VDD 802 810 VDD 796 VSS sky130_fd_sc_hd__or2_4 $T=162840 57120 1 0 $X=162650 $Y=54160
X2089 VSS VDD 836 618 VDD 829 VSS sky130_fd_sc_hd__or2_4 $T=165600 176800 0 0 $X=165410 $Y=176560
X2090 VSS VDD 885 875 VDD 879 VSS sky130_fd_sc_hd__or2_4 $T=176180 51680 0 0 $X=175990 $Y=51440
X2091 VSS VDD 899 851 VDD 893 VSS sky130_fd_sc_hd__or2_4 $T=177100 133280 0 0 $X=176910 $Y=133040
X2092 VSS VDD 867 912 VDD 886 VSS sky130_fd_sc_hd__or2_4 $T=177560 73440 1 0 $X=177370 $Y=70480
X2093 VSS VDD 920 830 VDD 807 VSS sky130_fd_sc_hd__or2_4 $T=183080 19040 0 0 $X=182890 $Y=18800
X2094 VSS VDD 774 848 VDD 934 VSS sky130_fd_sc_hd__or2_4 $T=189520 100640 1 0 $X=189330 $Y=97680
X2095 VSS VDD 963 912 VDD 959 VSS sky130_fd_sc_hd__or2_4 $T=193200 62560 1 0 $X=193010 $Y=59600
X2096 VSS VDD 1015 963 VDD 1008 VSS sky130_fd_sc_hd__or2_4 $T=205160 68000 1 0 $X=204970 $Y=65040
X2097 VSS VDD 1035 988 VDD 1015 VSS sky130_fd_sc_hd__or2_4 $T=209300 122400 1 0 $X=209110 $Y=119440
X2098 VSS VDD 997 973 VDD 1035 VSS sky130_fd_sc_hd__or2_4 $T=209300 138720 1 0 $X=209110 $Y=135760
X2099 VSS VDD 281 175 278 295 VDD 306 VSS sky130_fd_sc_hd__and4_4 $T=49220 127840 1 0 $X=49030 $Y=124880
X2100 VSS VDD 281 304 257 295 VDD 270 VSS sky130_fd_sc_hd__and4_4 $T=51520 133280 0 0 $X=51330 $Y=133040
X2101 VSS VDD 281 308 358 295 VDD 368 VSS sky130_fd_sc_hd__and4_4 $T=63020 127840 0 0 $X=62830 $Y=127600
X2102 VSS VDD 473 363 475 295 VDD 474 VSS sky130_fd_sc_hd__and4_4 $T=89240 138720 1 0 $X=89050 $Y=135760
X2103 VSS VDD 473 486 526 295 VDD 545 VSS sky130_fd_sc_hd__and4_4 $T=100280 144160 0 0 $X=100090 $Y=143920
X2104 VSS VDD 509 650 562 639 VDD 669 VSS sky130_fd_sc_hd__and4_4 $T=121900 89760 1 0 $X=121710 $Y=86800
X2105 VSS VDD 213 681 682 691 VDD 552 VSS sky130_fd_sc_hd__and4_4 $T=128800 193120 0 0 $X=128610 $Y=192880
X2106 VSS VDD 701 650 688 629 VDD 709 VSS sky130_fd_sc_hd__and4_4 $T=133400 73440 1 0 $X=133210 $Y=70480
X2107 VSS VDD 701 650 670 966 VDD 994 VSS sky130_fd_sc_hd__and4_4 $T=195040 51680 1 0 $X=194850 $Y=48720
X2108 VSS VDD 701 650 993 958 VDD 1018 VSS sky130_fd_sc_hd__and4_4 $T=201940 46240 1 0 $X=201750 $Y=43280
X2109 VSS VDD 701 985 1006 1008 VDD 1001 VSS sky130_fd_sc_hd__and4_4 $T=202860 73440 1 0 $X=202670 $Y=70480
X2110 VSS VDD 158 985 989 997 VDD 1021 VSS sky130_fd_sc_hd__and4_4 $T=202860 133280 1 0 $X=202670 $Y=130320
X2111 VSS VDD 701 985 1000 999 VDD 1027 VSS sky130_fd_sc_hd__and4_4 $T=203780 57120 1 0 $X=203590 $Y=54160
X2112 VSS VDD 158 985 1015 1022 VDD 1029 VSS sky130_fd_sc_hd__and4_4 $T=207920 116960 1 0 $X=207730 $Y=114000
X2113 VSS VDD 158 985 1039 1035 VDD 1030 VSS sky130_fd_sc_hd__and4_4 $T=208840 133280 0 0 $X=208650 $Y=133040
X2114 VSS VDD 279 298 238 ICV_32 $T=52900 19040 0 0 $X=52710 $Y=18800
X2115 VSS VDD 351 383 168 ICV_32 $T=66240 51680 1 0 $X=66050 $Y=48720
X2116 VSS VDD 355 388 SCAN_IN<18> ICV_32 $T=68080 116960 0 0 $X=67890 $Y=116720
X2117 VSS VDD 325 403 378 ICV_32 $T=69460 171360 0 0 $X=69270 $Y=171120
X2118 VSS VDD 371 420 437 ICV_32 $T=76820 214880 0 0 $X=76630 $Y=214640
X2119 VSS VDD 657 674 676 ICV_32 $T=124200 24480 0 0 $X=124010 $Y=24240
X2120 VSS VDD 801 337 836 ICV_32 $T=158700 176800 0 0 $X=158510 $Y=176560
X2121 VSS VDD 844 1046 1050 ICV_32 $T=208840 57120 1 0 $X=208650 $Y=54160
X2122 VSS VDD 68 39 68 39 VDD 75 VSS sky130_fd_sc_hd__a2bb2oi_4 $T=7820 160480 0 0 $X=7630 $Y=160240
X2123 VSS VDD 516 586 516 586 VDD 612 VSS sky130_fd_sc_hd__a2bb2oi_4 $T=111320 19040 1 0 $X=111130 $Y=16080
X2124 VSS VDD 981 974 981 974 VDD 1036 VSS sky130_fd_sc_hd__a2bb2oi_4 $T=206080 13600 0 0 $X=205890 $Y=13360
X2125 VSS VDD 995 996 995 996 VDD 1038 VSS sky130_fd_sc_hd__a2bb2oi_4 $T=208380 84320 0 0 $X=208190 $Y=84080
X2126 VSS VDD 1007 1017 1007 1017 VDD 1031 VSS sky130_fd_sc_hd__a2bb2oi_4 $T=208380 193120 0 0 $X=208190 $Y=192880
X2127 VSS VDD 44 ICV_33 $T=6900 78880 0 0 $X=6710 $Y=78640
X2128 VSS VDD 20 ICV_33 $T=14260 89760 0 0 $X=14070 $Y=89520
X2129 VSS VDD 96 ICV_33 $T=15180 176800 0 0 $X=14990 $Y=176560
X2130 VSS VDD 62 ICV_33 $T=16100 95200 0 0 $X=15910 $Y=94960
X2131 VSS VDD 104 ICV_33 $T=16100 182240 1 0 $X=15910 $Y=179280
X2132 VSS VDD SCAN_IN<10> ICV_33 $T=29440 116960 0 0 $X=29250 $Y=116720
X2133 VSS VDD 190 ICV_33 $T=29440 198560 1 0 $X=29250 $Y=195600
X2134 VSS VDD 179 ICV_33 $T=29900 78880 0 0 $X=29710 $Y=78640
X2135 VSS VDD 199 ICV_33 $T=30360 95200 1 0 $X=30170 $Y=92240
X2136 VSS VDD 203 ICV_33 $T=32660 24480 1 0 $X=32470 $Y=21520
X2137 VSS VDD 234 ICV_33 $T=38180 73440 0 0 $X=37990 $Y=73200
X2138 VSS VDD 275 ICV_33 $T=46000 62560 0 0 $X=45810 $Y=62320
X2139 VSS VDD 276 ICV_33 $T=46000 73440 0 0 $X=45810 $Y=73200
X2140 VSS VDD 257 ICV_33 $T=48300 133280 1 0 $X=48110 $Y=130320
X2141 VSS VDD 282 ICV_33 $T=48300 209440 1 0 $X=48110 $Y=206480
X2142 VSS VDD 84 ICV_33 $T=57960 29920 0 0 $X=57770 $Y=29680
X2143 VSS VDD 376 ICV_33 $T=66240 19040 1 0 $X=66050 $Y=16080
X2144 VSS VDD SCAN_IN<18> ICV_33 $T=73600 111520 0 0 $X=73410 $Y=111280
X2145 VSS VDD 413 ICV_33 $T=74520 133280 0 0 $X=74330 $Y=133040
X2146 VSS VDD 17 ICV_33 $T=82340 100640 0 0 $X=82150 $Y=100400
X2147 VSS VDD SCAN_IN<19> ICV_33 $T=86020 106080 0 0 $X=85830 $Y=105840
X2148 VSS VDD 17 ICV_33 $T=90160 62560 0 0 $X=89970 $Y=62320
X2149 VSS VDD 106 ICV_33 $T=91080 198560 1 0 $X=90890 $Y=195600
X2150 VSS VDD 501 ICV_33 $T=92920 46240 1 0 $X=92730 $Y=43280
X2151 VSS VDD 506 ICV_33 $T=95220 165920 0 0 $X=95030 $Y=165680
X2152 VSS VDD 17 ICV_33 $T=95680 29920 0 0 $X=95490 $Y=29680
X2153 VSS VDD 492 ICV_33 $T=100740 220320 0 0 $X=100550 $Y=220080
X2154 VSS VDD 550 ICV_33 $T=102120 176800 0 0 $X=101930 $Y=176560
X2155 VSS VDD 558 ICV_33 $T=103040 209440 0 0 $X=102850 $Y=209200
X2156 VSS VDD 565 ICV_33 $T=104420 73440 0 0 $X=104230 $Y=73200
X2157 VSS VDD 568 ICV_33 $T=104420 187680 0 0 $X=104230 $Y=187440
X2158 VSS VDD 591 ICV_33 $T=108100 57120 0 0 $X=107910 $Y=56880
X2159 VSS VDD 604 ICV_33 $T=113620 46240 0 0 $X=113430 $Y=46000
X2160 VSS VDD 20 ICV_33 $T=123280 122400 0 0 $X=123090 $Y=122160
X2161 VSS VDD 607 ICV_33 $T=124660 57120 0 0 $X=124470 $Y=56880
X2162 VSS VDD 213 ICV_33 $T=125120 193120 0 0 $X=124930 $Y=192880
X2163 VSS VDD 632 ICV_33 $T=126500 62560 1 0 $X=126310 $Y=59600
X2164 VSS VDD 674 ICV_33 $T=128340 29920 1 0 $X=128150 $Y=26960
X2165 VSS VDD 300 ICV_33 $T=128340 198560 0 0 $X=128150 $Y=198320
X2166 VSS VDD 671 ICV_33 $T=130180 220320 0 0 $X=129990 $Y=220080
X2167 VSS VDD 682 ICV_33 $T=132020 187680 0 0 $X=131830 $Y=187440
X2168 VSS VDD 487 ICV_33 $T=138920 84320 1 0 $X=138730 $Y=81360
X2169 VSS VDD 628 ICV_33 $T=142140 13600 0 0 $X=141950 $Y=13360
X2170 VSS VDD 764 ICV_33 $T=144440 13600 1 0 $X=144250 $Y=10640
X2171 VSS VDD 766 ICV_33 $T=149500 144160 1 0 $X=149310 $Y=141200
X2172 VSS VDD 608 ICV_33 $T=154560 89760 1 0 $X=154370 $Y=86800
X2173 VSS VDD 17 ICV_33 $T=154560 165920 0 0 $X=154370 $Y=165680
X2174 VSS VDD 792 ICV_33 $T=156400 171360 1 0 $X=156210 $Y=168400
X2175 VSS VDD 454 ICV_33 $T=157320 68000 0 0 $X=157130 $Y=67760
X2176 VSS VDD 834 ICV_33 $T=160540 182240 0 0 $X=160350 $Y=182000
X2177 VSS VDD 861 ICV_33 $T=170200 95200 0 0 $X=170010 $Y=94960
X2178 VSS VDD 851 ICV_33 $T=170200 127840 0 0 $X=170010 $Y=127600
X2179 VSS VDD 863 ICV_33 $T=174340 220320 1 0 $X=174150 $Y=217360
X2180 VSS VDD 887 ICV_33 $T=179400 51680 0 0 $X=179210 $Y=51440
X2181 VSS VDD 823 ICV_33 $T=184460 209440 1 0 $X=184270 $Y=206480
X2182 VSS VDD SCAN_IN<1> ICV_33 $T=185380 220320 0 0 $X=185190 $Y=220080
X2183 VSS VDD 801 ICV_33 $T=185840 182240 0 0 $X=185650 $Y=182000
X2184 VSS VDD SCAN_IN<5> ICV_33 $T=188600 165920 1 0 $X=188410 $Y=162960
X2185 VSS VDD 969 ICV_33 $T=194580 24480 0 0 $X=194390 $Y=24240
X2186 VSS VDD SCAN_IN<3> ICV_33 $T=195040 198560 0 0 $X=194850 $Y=198320
X2187 VSS VDD 963 ICV_33 $T=198260 68000 0 0 $X=198070 $Y=67760
X2188 VSS VDD 986 ICV_33 $T=198260 89760 0 0 $X=198070 $Y=89520
X2189 VSS VDD 1011 ICV_33 $T=201480 220320 1 0 $X=201290 $Y=217360
X2190 VSS VDD 981 ICV_33 $T=202400 13600 0 0 $X=202210 $Y=13360
X2191 VSS VDD 20 ICV_33 $T=202400 35360 0 0 $X=202210 $Y=35120
X2192 VSS VDD 979 ICV_33 $T=202400 193120 1 0 $X=202210 $Y=190160
X2193 VSS VDD 988 ICV_33 $T=207460 116960 0 0 $X=207270 $Y=116720
X2194 VSS VDD SCAN_IN<4> ICV_33 $T=208380 100640 0 0 $X=208190 $Y=100400
X2195 VSS VDD 10 21 20 VDD 84 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 29920 0 0 $X=7630 $Y=29680
X2196 VSS VDD 10 23 20 VDD 80 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 46240 0 0 $X=7630 $Y=46000
X2197 VSS VDD 10 45 20 VDD 98 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 116960 0 0 $X=7630 $Y=116720
X2198 VSS VDD CLK_OUT BB_IN RESET_N VDD DATA_OUT VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 122400 0 0 $X=7630 $Y=122160
X2199 VSS VDD 12 BB_IN RESET_N VDD 17 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 127840 0 0 $X=7630 $Y=127600
X2200 VSS VDD 14 46 RESET_N VDD 16 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 144160 0 0 $X=7630 $Y=143920
X2201 VSS VDD 17 18 RESET_N VDD 101 VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 214880 0 0 $X=7630 $Y=214640
X2202 VSS VDD 16 41 RESET_N VDD 110 VSS sky130_fd_sc_hd__dfrtp_4 $T=8740 220320 0 0 $X=8550 $Y=220080
X2203 VSS VDD 10 56 20 VDD 91 VSS sky130_fd_sc_hd__dfrtp_4 $T=9660 111520 0 0 $X=9470 $Y=111280
X2204 VSS VDD 10 71 20 VDD 129 VSS sky130_fd_sc_hd__dfrtp_4 $T=12420 68000 0 0 $X=12230 $Y=67760
X2205 VSS VDD 94 100 20 VDD 114 VSS sky130_fd_sc_hd__dfrtp_4 $T=17480 138720 0 0 $X=17290 $Y=138480
X2206 VSS VDD 10 86 20 VDD 172 VSS sky130_fd_sc_hd__dfrtp_4 $T=17940 89760 0 0 $X=17750 $Y=89520
X2207 VSS VDD 10 89 20 VDD 179 VSS sky130_fd_sc_hd__dfrtp_4 $T=19320 78880 0 0 $X=19130 $Y=78640
X2208 VSS VDD 10 178 20 VDD 251 VSS sky130_fd_sc_hd__dfrtp_4 $T=33580 35360 1 0 $X=33390 $Y=32400
X2209 VSS VDD 94 156 20 VDD 230 VSS sky130_fd_sc_hd__dfrtp_4 $T=34960 127840 0 0 $X=34770 $Y=127600
X2210 VSS VDD 10 185 20 VDD 261 VSS sky130_fd_sc_hd__dfrtp_4 $T=35420 46240 0 0 $X=35230 $Y=46000
X2211 VSS VDD 212 227 20 VDD 279 VSS sky130_fd_sc_hd__dfrtp_4 $T=38640 13600 0 0 $X=38450 $Y=13360
X2212 VSS VDD 94 270 20 VDD 324 VSS sky130_fd_sc_hd__dfrtp_4 $T=49220 138720 1 0 $X=49030 $Y=135760
X2213 VSS VDD 94 293 20 VDD 272 VSS sky130_fd_sc_hd__dfrtp_4 $T=49220 176800 1 0 $X=49030 $Y=173840
X2214 VSS VDD 212 17 20 VDD 334 VSS sky130_fd_sc_hd__dfrtp_4 $T=51520 106080 1 0 $X=51330 $Y=103120
X2215 VSS VDD 94 306 20 VDD 355 VSS sky130_fd_sc_hd__dfrtp_4 $T=53820 122400 1 0 $X=53630 $Y=119440
X2216 VSS VDD 212 169 20 VDD 365 VSS sky130_fd_sc_hd__dfrtp_4 $T=55660 19040 1 0 $X=55470 $Y=16080
X2217 VSS VDD 212 352 20 VDD CLK_OUT VSS sky130_fd_sc_hd__dfrtp_4 $T=63020 111520 0 0 $X=62830 $Y=111280
X2218 VSS VDD 94 368 20 VDD 388 VSS sky130_fd_sc_hd__dfrtp_4 $T=64400 122400 0 0 $X=64210 $Y=122160
X2219 VSS VDD 212 393 20 VDD 421 VSS sky130_fd_sc_hd__dfrtp_4 $T=70840 89760 0 0 $X=70650 $Y=89520
X2220 VSS VDD 94 474 20 VDD 377 VSS sky130_fd_sc_hd__dfrtp_4 $T=89700 122400 1 0 $X=89510 $Y=119440
X2221 VSS VDD 456 468 20 VDD 460 VSS sky130_fd_sc_hd__dfrtp_4 $T=91080 155040 0 0 $X=90890 $Y=154800
X2222 VSS VDD 456 567 20 VDD 607 VSS sky130_fd_sc_hd__dfrtp_4 $T=105340 100640 1 0 $X=105150 $Y=97680
X2223 VSS VDD 456 569 20 VDD 558 VSS sky130_fd_sc_hd__dfrtp_4 $T=105340 160480 1 0 $X=105150 $Y=157520
X2224 VSS VDD 456 545 20 VDD 618 VSS sky130_fd_sc_hd__dfrtp_4 $T=108560 144160 1 0 $X=108370 $Y=141200
X2225 VSS VDD 456 662 20 VDD 673 VSS sky130_fd_sc_hd__dfrtp_4 $T=123740 144160 0 0 $X=123550 $Y=143920
X2226 VSS VDD 456 667 20 VDD 678 VSS sky130_fd_sc_hd__dfrtp_4 $T=124660 160480 0 0 $X=124470 $Y=160240
X2227 VSS VDD 456 669 20 VDD 672 VSS sky130_fd_sc_hd__dfrtp_4 $T=126500 89760 0 0 $X=126310 $Y=89520
X2228 VSS VDD 416 659 20 VDD 723 VSS sky130_fd_sc_hd__dfrtp_4 $T=126960 122400 0 0 $X=126770 $Y=122160
X2229 VSS VDD 456 689 20 VDD 731 VSS sky130_fd_sc_hd__dfrtp_4 $T=130180 78880 0 0 $X=129990 $Y=78640
X2230 VSS VDD 456 709 20 VDD 666 VSS sky130_fd_sc_hd__dfrtp_4 $T=133400 78880 1 0 $X=133210 $Y=75920
X2231 VSS VDD 16 495 20 VDD 747 VSS sky130_fd_sc_hd__dfrtp_4 $T=145820 220320 1 0 $X=145630 $Y=217360
X2232 VSS VDD 16 683 20 VDD 795 VSS sky130_fd_sc_hd__dfrtp_4 $T=154100 214880 0 0 $X=153910 $Y=214640
X2233 VSS VDD 17 871 20 VDD 929 VSS sky130_fd_sc_hd__dfrtp_4 $T=173880 160480 1 0 $X=173690 $Y=157520
X2234 VSS VDD 17 870 20 VDD 960 VSS sky130_fd_sc_hd__dfrtp_4 $T=182160 160480 0 0 $X=181970 $Y=160240
X2235 VSS VDD 844 994 20 VDD 904 VSS sky130_fd_sc_hd__dfrtp_4 $T=203320 46240 0 0 $X=203130 $Y=46000
X2236 VSS VDD 844 1001 20 VDD 987 VSS sky130_fd_sc_hd__dfrtp_4 $T=203780 73440 0 0 $X=203590 $Y=73200
X2237 VSS VDD 844 1021 20 VDD 940 VSS sky130_fd_sc_hd__dfrtp_4 $T=205620 127840 0 0 $X=205430 $Y=127600
X2238 VSS VDD 844 1018 20 VDD 765 VSS sky130_fd_sc_hd__dfrtp_4 $T=206080 35360 0 0 $X=205890 $Y=35120
X2239 VSS VDD 844 1027 20 VDD 911 VSS sky130_fd_sc_hd__dfrtp_4 $T=207460 51680 0 0 $X=207270 $Y=51440
X2240 VSS VDD 844 1029 20 VDD 977 VSS sky130_fd_sc_hd__dfrtp_4 $T=207460 111520 0 0 $X=207270 $Y=111280
X2241 VSS VDD 844 1030 20 VDD 1003 VSS sky130_fd_sc_hd__dfrtp_4 $T=207460 122400 0 0 $X=207270 $Y=122160
X2242 VSS VDD 73 119 88 54 ICV_34 $T=19320 46240 0 0 $X=19130 $Y=46000
X2243 VSS VDD 159 120 159 155 ICV_34 $T=26220 116960 1 0 $X=26030 $Y=114000
X2244 VSS VDD 106 547 106 540 ICV_34 $T=104420 193120 0 0 $X=104230 $Y=192880
X2245 VSS VDD 558 558 460 549 ICV_34 $T=106720 160480 0 0 $X=106530 $Y=160240
X2246 VSS VDD 625 673 625 561 ICV_34 $T=125120 149600 0 0 $X=124930 $Y=149360
X2247 VSS VDD 641 738 680 653 ICV_34 $T=139380 187680 1 0 $X=139190 $Y=184720
X2248 VSS VDD 747 747 770 696 ICV_34 $T=151340 204000 0 0 $X=151150 $Y=203760
X2249 VSS VDD 756 865 756 897 ICV_34 $T=174340 35360 1 0 $X=174150 $Y=32400
X2250 VSS VDD 1027 911 1037 1041 ICV_34 $T=207460 51680 1 0 $X=207270 $Y=48720
X2251 VSS 59 87 143 ICV_35 $T=22080 187680 1 0 $X=21890 $Y=184720
X2252 VSS 266 211 242 ICV_35 $T=41860 89760 0 0 $X=41670 $Y=89520
X2253 VSS 55 267 216 ICV_35 $T=51520 84320 1 0 $X=51330 $Y=81360
X2254 VSS 290 343 349 ICV_35 $T=63020 214880 0 0 $X=62830 $Y=214640
X2255 VSS 20 507 456 ICV_35 $T=119140 160480 0 0 $X=118950 $Y=160240
X2256 VSS 902 911 958 ICV_35 $T=188600 46240 0 0 $X=188410 $Y=46000
X2257 VSS 973 989 985 ICV_35 $T=203320 133280 0 0 $X=203130 $Y=133040
X2258 VSS 911 930 999 ICV_35 $T=207460 40800 0 0 $X=207270 $Y=40560
X2259 VSS VDD 122 103 90 95 VDD 104 VSS sky130_fd_sc_hd__a211o_4 $T=18860 165920 0 0 $X=18670 $Y=165680
X2260 VSS VDD 180 155 177 152 VDD 140 VSS sky130_fd_sc_hd__a211o_4 $T=26680 111520 1 0 $X=26490 $Y=108560
X2261 VSS VDD 114 174 118 173 VDD 184 VSS sky130_fd_sc_hd__a211o_4 $T=31280 165920 1 0 $X=31090 $Y=162960
X2262 VSS VDD 201 140 194 91 VDD 205 VSS sky130_fd_sc_hd__a211o_4 $T=34960 100640 0 0 $X=34770 $Y=100400
X2263 VSS VDD 210 192 181 43 VDD 224 VSS sky130_fd_sc_hd__a211o_4 $T=37720 68000 1 0 $X=37530 $Y=65040
X2264 VSS VDD 239 254 223 265 VDD 288 VSS sky130_fd_sc_hd__a211o_4 $T=49680 57120 1 0 $X=49490 $Y=54160
X2265 VSS VDD 298 287 288 274 VDD 260 VSS sky130_fd_sc_hd__a211o_4 $T=51520 24480 0 0 $X=51330 $Y=24240
X2266 VSS VDD 298 317 238 191 VDD 322 VSS sky130_fd_sc_hd__a211o_4 $T=57960 24480 1 0 $X=57770 $Y=21520
X2267 VSS VDD 84 191 361 251 VDD 332 VSS sky130_fd_sc_hd__a211o_4 $T=60260 35360 1 0 $X=60070 $Y=32400
X2268 VSS VDD 333 318 351 307 VDD 273 VSS sky130_fd_sc_hd__a211o_4 $T=63020 51680 0 0 $X=62830 $Y=51440
X2269 VSS VDD 392 387 168 373 VDD 366 VSS sky130_fd_sc_hd__a211o_4 $T=69000 62560 0 0 $X=68810 $Y=62320
X2270 VSS VDD 385 394 378 349 VDD 395 VSS sky130_fd_sc_hd__a211o_4 $T=71300 187680 0 0 $X=71110 $Y=187440
X2271 VSS VDD 438 439 356 422 VDD 431 VSS sky130_fd_sc_hd__a211o_4 $T=79580 122400 1 0 $X=79390 $Y=119440
X2272 VSS VDD 237 419 580 552 VDD 222 VSS sky130_fd_sc_hd__a211o_4 $T=105340 187680 1 0 $X=105150 $Y=184720
X2273 VSS VDD 603 611 570 573 VDD 577 VSS sky130_fd_sc_hd__a211o_4 $T=113620 29920 1 0 $X=113430 $Y=26960
X2274 VSS VDD 615 575 618 644 VDD 478 VSS sky130_fd_sc_hd__a211o_4 $T=116840 122400 1 0 $X=116650 $Y=119440
X2275 VSS VDD 485 555 624 SCAN_IN<14> VDD 594 VSS sky130_fd_sc_hd__a211o_4 $T=119140 133280 0 0 $X=118950 $Y=133040
X2276 VSS VDD 651 640 568 547 VDD 619 VSS sky130_fd_sc_hd__a211o_4 $T=121900 182240 1 0 $X=121710 $Y=179280
X2277 VSS VDD 607 687 632 534 VDD 677 VSS sky130_fd_sc_hd__a211o_4 $T=128340 57120 0 0 $X=128150 $Y=56880
X2278 VSS VDD 653 715 624 690 VDD 686 VSS sky130_fd_sc_hd__a211o_4 $T=134780 182240 0 0 $X=134590 $Y=182000
X2279 VSS VDD 739 705 733 721 VDD 722 VSS sky130_fd_sc_hd__a211o_4 $T=136160 133280 1 0 $X=135970 $Y=130320
X2280 VSS VDD 768 726 422 756 VDD 702 VSS sky130_fd_sc_hd__a211o_4 $T=147200 95200 0 0 $X=147010 $Y=94960
X2281 VSS VDD 743 772 758 757 VDD 732 VSS sky130_fd_sc_hd__a211o_4 $T=147200 122400 0 0 $X=147010 $Y=122160
X2282 VSS VDD 901 868 877 558 VDD 889 VSS sky130_fd_sc_hd__a211o_4 $T=171580 214880 1 0 $X=171390 $Y=211920
X2283 VSS VDD 1012 1016 1044 940 VDD 1025 VSS sky130_fd_sc_hd__a211o_4 $T=207000 171360 0 0 $X=206810 $Y=171120
X2284 VSS VDD 11 ICV_36 $T=6900 89760 0 0 $X=6710 $Y=89520
X2285 VSS VDD 57 ICV_36 $T=10580 176800 0 0 $X=10390 $Y=176560
X2286 VSS VDD 20 ICV_36 $T=14260 138720 0 0 $X=14070 $Y=138480
X2287 VSS VDD 105 ICV_36 $T=18860 182240 0 0 $X=18670 $Y=182000
X2288 VSS VDD 155 ICV_36 $T=23920 106080 1 0 $X=23730 $Y=103120
X2289 VSS VDD 102 ICV_36 $T=31740 182240 1 0 $X=31550 $Y=179280
X2290 VSS VDD 201 ICV_36 $T=32660 106080 1 0 $X=32470 $Y=103120
X2291 VSS VDD 149 ICV_36 $T=34040 182240 0 0 $X=33850 $Y=182000
X2292 VSS VDD 181 ICV_36 $T=36340 62560 1 0 $X=36150 $Y=59600
X2293 VSS VDD 285 ICV_36 $T=48300 106080 1 0 $X=48110 $Y=103120
X2294 VSS VDD 308 ICV_36 $T=51520 127840 0 0 $X=51330 $Y=127600
X2295 VSS VDD 315 ICV_36 $T=53360 127840 1 0 $X=53170 $Y=124880
X2296 VSS VDD 26 ICV_36 $T=55200 78880 1 0 $X=55010 $Y=75920
X2297 VSS VDD 324 ICV_36 $T=56120 138720 0 0 $X=55930 $Y=138480
X2298 VSS VDD 251 ICV_36 $T=62100 35360 0 0 $X=61910 $Y=35120
X2299 VSS VDD 347 ICV_36 $T=62100 138720 0 0 $X=61910 $Y=138480
X2300 VSS VDD 324 ICV_36 $T=62100 165920 0 0 $X=61910 $Y=165680
X2301 VSS VDD 330 ICV_36 $T=65780 57120 0 0 $X=65590 $Y=56880
X2302 VSS VDD 20 ICV_36 $T=67620 89760 0 0 $X=67430 $Y=89520
X2303 VSS VDD 380 ICV_36 $T=67620 106080 1 0 $X=67430 $Y=103120
X2304 VSS VDD 385 ICV_36 $T=68080 187680 0 0 $X=67890 $Y=187440
X2305 VSS VDD 370 ICV_36 $T=69920 106080 1 0 $X=69730 $Y=103120
X2306 VSS VDD 441 ICV_36 $T=86480 165920 0 0 $X=86290 $Y=165680
X2307 VSS VDD 470 ICV_36 $T=86480 198560 0 0 $X=86290 $Y=198320
X2308 VSS VDD 513 ICV_36 $T=95680 46240 0 0 $X=95490 $Y=46000
X2309 VSS VDD 417 ICV_36 $T=95680 73440 0 0 $X=95490 $Y=73200
X2310 VSS VDD 514 ICV_36 $T=96140 24480 1 0 $X=95950 $Y=21520
X2311 VSS VDD 50 ICV_36 $T=100280 19040 1 0 $X=100090 $Y=16080
X2312 VSS VDD 534 ICV_36 $T=100280 62560 1 0 $X=100090 $Y=59600
X2313 VSS VDD 588 ICV_36 $T=108100 106080 1 0 $X=107910 $Y=103120
X2314 VSS VDD 607 ICV_36 $T=112240 73440 0 0 $X=112050 $Y=73200
X2315 VSS VDD 619 ICV_36 $T=114540 182240 0 0 $X=114350 $Y=182000
X2316 VSS VDD 648 ICV_36 $T=120060 100640 0 0 $X=119870 $Y=100400
X2317 VSS VDD 635 ICV_36 $T=122820 176800 0 0 $X=122630 $Y=176560
X2318 VSS VDD 713 ICV_36 $T=132940 204000 0 0 $X=132750 $Y=203760
X2319 VSS VDD 622 ICV_36 $T=138920 51680 0 0 $X=138730 $Y=51440
X2320 VSS VDD 741 ICV_36 $T=141220 165920 1 0 $X=141030 $Y=162960
X2321 VSS VDD 758 ICV_36 $T=144900 127840 1 0 $X=144710 $Y=124880
X2322 VSS VDD 16 ICV_36 $T=146280 182240 0 0 $X=146090 $Y=182000
X2323 VSS VDD 756 ICV_36 $T=148120 68000 0 0 $X=147930 $Y=67760
X2324 VSS VDD 520 ICV_36 $T=150420 78880 0 0 $X=150230 $Y=78640
X2325 VSS VDD 791 ICV_36 $T=153180 149600 0 0 $X=152990 $Y=149360
X2326 VSS VDD 745 ICV_36 $T=156400 116960 1 0 $X=156210 $Y=114000
X2327 VSS VDD 568 ICV_36 $T=156860 176800 1 0 $X=156670 $Y=173840
X2328 VSS VDD 814 ICV_36 $T=160540 155040 1 0 $X=160350 $Y=152080
X2329 VSS VDD 802 ICV_36 $T=164680 73440 1 0 $X=164490 $Y=70480
X2330 VSS VDD 532 ICV_36 $T=168820 171360 0 0 $X=168630 $Y=171120
X2331 VSS VDD 20 ICV_36 $T=180780 165920 1 0 $X=180590 $Y=162960
X2332 VSS VDD 721 ICV_36 $T=182160 138720 0 0 $X=181970 $Y=138480
X2333 VSS VDD 771 ICV_36 $T=182620 62560 0 0 $X=182430 $Y=62320
X2334 VSS VDD 942 ICV_36 $T=184460 133280 1 0 $X=184270 $Y=130320
X2335 VSS VDD SCAN_IN<3> ICV_36 $T=187220 193120 0 0 $X=187030 $Y=192880
X2336 VSS VDD 972 ICV_36 $T=192280 116960 1 0 $X=192090 $Y=114000
X2337 VSS VDD 920 ICV_36 $T=195040 13600 1 0 $X=194850 $Y=10640
X2338 VSS VDD 1006 ICV_36 $T=199640 73440 1 0 $X=199450 $Y=70480
X2339 VSS VDD 1004 ICV_36 $T=202400 19040 0 0 $X=202210 $Y=18800
X2340 VSS VDD 20 ICV_36 $T=202400 127840 0 0 $X=202210 $Y=127600
X2341 VSS VDD 765 ICV_36 $T=206080 29920 0 0 $X=205890 $Y=29680
X2342 VSS VDD 1030 ICV_36 $T=206080 122400 1 0 $X=205890 $Y=119440
X2343 VSS VDD 1014 ICV_36 $T=206080 198560 0 0 $X=205890 $Y=198320
X2344 VSS VDD 973 ICV_36 $T=207000 138720 0 0 $X=206810 $Y=138480
X2345 VSS VDD 19 ICV_37 $T=7820 24480 1 0 $X=7630 $Y=21520
X2346 VSS VDD 24 ICV_37 $T=7820 62560 1 0 $X=7630 $Y=59600
X2347 VSS VDD 24 ICV_37 $T=7820 73440 1 0 $X=7630 $Y=70480
X2348 VSS VDD 20 ICV_37 $T=7820 187680 1 0 $X=7630 $Y=184720
X2349 VSS VDD 11 ICV_37 $T=12880 100640 0 0 $X=12690 $Y=100400
X2350 VSS VDD 84 ICV_37 $T=14720 24480 0 0 $X=14530 $Y=24240
X2351 VSS VDD 100 ICV_37 $T=17480 144160 1 0 $X=17290 $Y=141200
X2352 VSS VDD 88 ICV_37 $T=21160 46240 1 0 $X=20970 $Y=43280
X2353 VSS VDD 122 ICV_37 $T=21160 171360 1 0 $X=20970 $Y=168400
X2354 VSS VDD 114 ICV_37 $T=31280 160480 0 0 $X=31090 $Y=160240
X2355 VSS VDD 95 ICV_37 $T=37260 144160 0 0 $X=37070 $Y=143920
X2356 VSS VDD 285 ICV_37 $T=59340 78880 0 0 $X=59150 $Y=78640
X2357 VSS VDD 343 ICV_37 $T=62100 225760 1 0 $X=61910 $Y=222800
X2358 VSS VDD 332 ICV_37 $T=63020 62560 0 0 $X=62830 $Y=62320
X2359 VSS VDD 330 ICV_37 $T=63020 73440 0 0 $X=62830 $Y=73200
X2360 VSS VDD 366 ICV_37 $T=66700 68000 1 0 $X=66510 $Y=65040
X2361 VSS VDD 150 ICV_37 $T=74060 198560 0 0 $X=73870 $Y=198320
X2362 VSS VDD 414 ICV_37 $T=76360 171360 0 0 $X=76170 $Y=171120
X2363 VSS VDD 422 ICV_37 $T=77280 116960 1 0 $X=77090 $Y=114000
X2364 VSS VDD 315 ICV_37 $T=77280 122400 1 0 $X=77090 $Y=119440
X2365 VSS VDD 357 ICV_37 $T=87400 209440 0 0 $X=87210 $Y=209200
X2366 VSS VDD 464 ICV_37 $T=87400 220320 0 0 $X=87210 $Y=220080
X2367 VSS VDD 533 ICV_37 $T=101660 24480 1 0 $X=101470 $Y=21520
X2368 VSS VDD 517 ICV_37 $T=101660 133280 1 0 $X=101470 $Y=130320
X2369 VSS VDD 401 ICV_37 $T=101660 198560 1 0 $X=101470 $Y=195600
X2370 VSS VDD 145 ICV_37 $T=101660 204000 1 0 $X=101470 $Y=201040
X2371 VSS VDD 559 ICV_37 $T=105340 68000 1 0 $X=105150 $Y=65040
X2372 VSS VDD 491 ICV_37 $T=109480 204000 1 0 $X=109290 $Y=201040
X2373 VSS VDD 591 ICV_37 $T=110860 68000 1 0 $X=110670 $Y=65040
X2374 VSS VDD 58 ICV_37 $T=115460 198560 0 0 $X=115270 $Y=198320
X2375 VSS VDD 547 ICV_37 $T=123740 176800 1 0 $X=123550 $Y=173840
X2376 VSS VDD 633 ICV_37 $T=133400 187680 1 0 $X=133210 $Y=184720
X2377 VSS VDD 736 ICV_37 $T=143520 89760 0 0 $X=143330 $Y=89520
X2378 VSS VDD 464 ICV_37 $T=143520 220320 1 0 $X=143330 $Y=217360
X2379 VSS VDD 738 ICV_37 $T=146280 198560 1 0 $X=146090 $Y=195600
X2380 VSS VDD 620 ICV_37 $T=147200 187680 0 0 $X=147010 $Y=187440
X2381 VSS VDD 551 ICV_37 $T=157780 122400 1 0 $X=157590 $Y=119440
X2382 VSS VDD 886 ICV_37 $T=175260 68000 0 0 $X=175070 $Y=67760
X2383 VSS VDD 905 ICV_37 $T=177100 182240 1 0 $X=176910 $Y=179280
X2384 VSS VDD 947 ICV_37 $T=193200 193120 0 0 $X=193010 $Y=192880
X2385 VSS VDD 960 ICV_37 $T=196880 155040 1 0 $X=196690 $Y=152080
X2386 VSS VDD 930 ICV_37 $T=203780 35360 1 0 $X=203590 $Y=32400
X2387 VSS VDD 940 ICV_37 $T=205620 155040 0 0 $X=205430 $Y=154800
X2388 VSS VDD 981 ICV_37 $T=206080 19040 1 0 $X=205890 $Y=16080
X2389 VSS VDD 844 ICV_37 $T=207000 46240 1 0 $X=206810 $Y=43280
X2390 VSS VDD 24 19 ICV_38 $T=8280 57120 1 0 $X=8090 $Y=54160
X2391 VSS VDD 160 113 ICV_38 $T=26680 127840 1 0 $X=26490 $Y=124880
X2392 VSS VDD 279 191 ICV_38 $T=49680 19040 1 0 $X=49490 $Y=16080
X2393 VSS VDD 272 92 ICV_38 $T=52440 209440 1 0 $X=52250 $Y=206480
X2394 VSS VDD 307 168 ICV_38 $T=55200 46240 1 0 $X=55010 $Y=43280
X2395 VSS VDD 325 349 ICV_38 $T=66700 176800 1 0 $X=66510 $Y=173840
X2396 VSS VDD 357 321 ICV_38 $T=81420 209440 1 0 $X=81230 $Y=206480
X2397 VSS VDD 17 448 ICV_38 $T=93380 73440 1 0 $X=93190 $Y=70480
X2398 VSS VDD 678 507 ICV_38 $T=136160 165920 1 0 $X=135970 $Y=162960
X2399 VSS VDD 855 633 ICV_38 $T=166520 225760 1 0 $X=166330 $Y=222800
X2400 VSS VDD 976 848 ICV_38 $T=195500 100640 1 0 $X=195310 $Y=97680
X2401 VSS VDD 977 776 ICV_38 $T=195500 111520 1 0 $X=195310 $Y=108560
X2402 VSS VDD 969 875 ICV_38 $T=198260 35360 1 0 $X=198070 $Y=32400
X2403 VSS VDD 1024 930 ICV_38 $T=207000 29920 1 0 $X=206810 $Y=26960
X2404 VSS RESET_N 46 67 82 ICV_39 $T=7820 149600 1 0 $X=7630 $Y=146640
X2405 VSS 31 57 50 50 ICV_39 $T=7820 155040 1 0 $X=7630 $Y=152080
X2406 VSS 36 37 64 62 ICV_39 $T=8280 84320 0 0 $X=8090 $Y=84080
X2407 VSS SCAN_IN<9> 33 69 68 ICV_39 $T=8740 165920 1 0 $X=8550 $Y=162960
X2408 VSS 59 76 83 92 ICV_39 $T=10120 187680 1 0 $X=9930 $Y=184720
X2409 VSS 39 118 131 75 ICV_39 $T=18400 160480 0 0 $X=18210 $Y=160240
X2410 VSS 112 120 64 37 ICV_39 $T=19320 84320 0 0 $X=19130 $Y=84080
X2411 VSS 130 SCAN_IN<10> 105 173 ICV_39 $T=22080 144160 0 0 $X=21890 $Y=143920
X2412 VSS 144 59 150 166 ICV_39 $T=23920 193120 0 0 $X=23730 $Y=192880
X2413 VSS 109 175 158 20 ICV_39 $T=26220 127840 0 0 $X=26030 $Y=127600
X2414 VSS 60 198 119 210 ICV_39 $T=30360 68000 1 0 $X=30170 $Y=65040
X2415 VSS 189 118 127 118 ICV_39 $T=31280 193120 1 0 $X=31090 $Y=190160
X2416 VSS 180 217 194 214 ICV_39 $T=34960 106080 0 0 $X=34770 $Y=105840
X2417 VSS 254 265 273 239 ICV_39 $T=43700 51680 0 0 $X=43510 $Y=51440
X2418 VSS 295 175 299 308 ICV_39 $T=51520 122400 0 0 $X=51330 $Y=122160
X2419 VSS 252 292 319 329 ICV_39 $T=52440 155040 0 0 $X=52250 $Y=154800
X2420 VSS 37 266 266 37 ICV_39 $T=53820 84320 0 0 $X=53630 $Y=84080
X2421 VSS 314 321 166 340 ICV_39 $T=54280 198560 0 0 $X=54090 $Y=198320
X2422 VSS 347 363 355 377 ICV_39 $T=63020 133280 0 0 $X=62830 $Y=133040
X2423 VSS 374 349 396 399 ICV_39 $T=67160 214880 1 0 $X=66970 $Y=211920
X2424 VSS 409 114 230 404 ICV_39 $T=74520 138720 0 0 $X=74330 $Y=138480
X2425 VSS 410 339 364 378 ICV_39 $T=74520 165920 0 0 $X=74330 $Y=165680
X2426 VSS 412 365 386 147 ICV_39 $T=76360 19040 0 0 $X=76170 $Y=18800
X2427 VSS 213 300 426 446 ICV_39 $T=78660 187680 0 0 $X=78470 $Y=187440
X2428 VSS 432 188 230 449 ICV_39 $T=79120 127840 0 0 $X=78930 $Y=127600
X2429 VSS 536 548 346 565 ICV_39 $T=102120 89760 0 0 $X=101930 $Y=89520
X2430 VSS 419 552 237 580 ICV_39 $T=102580 182240 0 0 $X=102390 $Y=182000
X2431 VSS 544 553 401 581 ICV_39 $T=102580 214880 0 0 $X=102390 $Y=214640
X2432 VSS 512 SCAN_IN<15> 377 589 ICV_39 $T=103960 116960 0 0 $X=103770 $Y=116720
X2433 VSS 537 494 517 594 ICV_39 $T=105340 127840 0 0 $X=105150 $Y=127600
X2434 VSS 551 587 593 564 ICV_39 $T=107180 35360 0 0 $X=106990 $Y=35120
X2435 VSS 547 557 515 401 ICV_39 $T=108100 198560 0 0 $X=107910 $Y=198320
X2436 VSS 20 545 456 476 ICV_39 $T=108560 138720 0 0 $X=108370 $Y=138480
X2437 VSS 633 634 595 290 ICV_39 $T=119140 214880 0 0 $X=118950 $Y=214640
X2438 VSS 636 489 623 668 ICV_39 $T=120060 35360 0 0 $X=119870 $Y=35120
X2439 VSS 679 253 676 SCAN_IN<8> ICV_39 $T=128800 13600 0 0 $X=128610 $Y=13360
X2440 VSS 680 693 SCAN_IN<13> 673 ICV_39 $T=128800 138720 0 0 $X=128610 $Y=138480
X2441 VSS 648 664 710 702 ICV_39 $T=130640 100640 0 0 $X=130450 $Y=100400
X2442 VSS 637 650 701 629 ICV_39 $T=132020 68000 0 0 $X=131830 $Y=67760
X2443 VSS 672 449 717 711 ICV_39 $T=133860 106080 0 0 $X=133670 $Y=105840
X2444 VSS 712 346 728 734 ICV_39 $T=134320 149600 0 0 $X=134130 $Y=149360
X2445 VSS 720 732 743 753 ICV_39 $T=137080 116960 0 0 $X=136890 $Y=116720
X2446 VSS 741 750 507 761 ICV_39 $T=144440 171360 1 0 $X=144250 $Y=168400
X2447 VSS 772 737 776 693 ICV_39 $T=147200 116960 0 0 $X=147010 $Y=116720
X2448 VSS 781 698 574 805 ICV_39 $T=151340 40800 1 0 $X=151150 $Y=37840
X2449 VSS 806 812 698 832 ICV_39 $T=156860 95200 0 0 $X=156670 $Y=94960
X2450 VSS 596 831 698 850 ICV_39 $T=160540 73440 0 0 $X=160350 $Y=73200
X2451 VSS 787 703 849 858 ICV_39 $T=161460 111520 1 0 $X=161270 $Y=108560
X2452 VSS 788 756 830 810 ICV_39 $T=161920 29920 0 0 $X=161730 $Y=29680
X2453 VSS 828 839 852 790 ICV_39 $T=161920 149600 1 0 $X=161730 $Y=146640
X2454 VSS 857 873 624 20 ICV_39 $T=166520 193120 0 0 $X=166330 $Y=192880
X2455 VSS 898 848 17 20 ICV_39 $T=172500 100640 1 0 $X=172310 $Y=97680
X2456 VSS 865 830 880 17 ICV_39 $T=176180 24480 0 0 $X=175990 $Y=24240
X2457 VSS 939 943 757 851 ICV_39 $T=184920 133280 0 0 $X=184730 $Y=133040
X2458 VSS 875 930 954 962 ICV_39 $T=189060 35360 0 0 $X=188870 $Y=35120
X2459 VSS 760 953 953 935 ICV_39 $T=193660 19040 0 0 $X=193470 $Y=18800
X2460 VSS 971 927 988 982 ICV_39 $T=193660 111520 0 0 $X=193470 $Y=111280
X2461 VSS 975 913 973 983 ICV_39 $T=194120 138720 0 0 $X=193930 $Y=138480
X2462 VSS 917 SCAN_IN<1> 819 915 ICV_39 $T=194120 176800 0 0 $X=193930 $Y=176560
X2463 VSS 923 967 927 977 ICV_39 $T=194580 116960 0 0 $X=194390 $Y=116720
X2464 VSS 1002 914 986 976 ICV_39 $T=200100 95200 1 0 $X=199910 $Y=92240
X2465 VSS 1017 1017 1007 1026 ICV_39 $T=204700 198560 1 0 $X=204510 $Y=195600
X2466 VSS 974 1024 974 1036 ICV_39 $T=206540 13600 1 0 $X=206350 $Y=10640
X2467 VSS VDD 10 28 56 ICV_40 $T=7820 111520 1 0 $X=7630 $Y=108560
X2468 VSS VDD 10 20 45 ICV_40 $T=7820 116960 1 0 $X=7630 $Y=114000
X2469 VSS VDD RESET_N BB_IN CLK_OUT ICV_40 $T=7820 122400 1 0 $X=7630 $Y=119440
X2470 VSS VDD 18 RESET_N 17 ICV_40 $T=7820 214880 1 0 $X=7630 $Y=211920
X2471 VSS VDD 166 125 150 ICV_40 $T=23000 187680 0 0 $X=22810 $Y=187440
X2472 VSS VDD 117 168 157 ICV_40 $T=30360 40800 1 0 $X=30170 $Y=37840
X2473 VSS VDD 246 204 210 ICV_40 $T=39100 57120 0 0 $X=38910 $Y=56880
X2474 VSS VDD 212 214 20 ICV_40 $T=49680 100640 1 0 $X=49490 $Y=97680
X2475 VSS VDD 212 20 296 ICV_40 $T=49680 106080 0 0 $X=49490 $Y=105840
X2476 VSS VDD 280 145 305 ICV_40 $T=50140 214880 0 0 $X=49950 $Y=214640
X2477 VSS VDD 94 20 281 ICV_40 $T=64400 127840 1 0 $X=64210 $Y=124880
X2478 VSS VDD 411 16 20 ICV_40 $T=76360 198560 0 0 $X=76170 $Y=198320
X2479 VSS VDD 92 415 301 ICV_40 $T=76360 209440 0 0 $X=76170 $Y=209200
X2480 VSS VDD 429 418 407 ICV_40 $T=77280 160480 1 0 $X=77090 $Y=157520
X2481 VSS VDD 395 385 389 ICV_40 $T=77280 182240 0 0 $X=77090 $Y=182000
X2482 VSS VDD 416 20 440 ICV_40 $T=79580 62560 0 0 $X=79390 $Y=62320
X2483 VSS VDD 479 476 482 ICV_40 $T=89700 160480 1 0 $X=89510 $Y=157520
X2484 VSS VDD 485 486 476 ICV_40 $T=92460 138720 0 0 $X=92270 $Y=138480
X2485 VSS VDD 433 499 481 ICV_40 $T=93840 171360 0 0 $X=93650 $Y=171120
X2486 VSS VDD 245 357 240 ICV_40 $T=105340 209440 1 0 $X=105150 $Y=206480
X2487 VSS VDD 649 707 695 ICV_40 $T=133860 46240 0 0 $X=133670 $Y=46000
X2488 VSS VDD 774 771 774 ICV_40 $T=147200 106080 1 0 $X=147010 $Y=103120
X2489 VSS VDD 690 20 601 ICV_40 $T=149500 182240 1 0 $X=149310 $Y=179280
X2490 VSS VDD 963 875 959 ICV_40 $T=189520 57120 1 0 $X=189330 $Y=54160
X2491 VSS VDD 964 912 963 ICV_40 $T=190900 62560 0 0 $X=190710 $Y=62320
X2492 VSS VDD 844 1021 844 ICV_40 $T=205620 127840 1 0 $X=205430 $Y=124880
X2493 VSS VDD 1012 SCAN_IN<1> 819 ICV_40 $T=206080 176800 0 0 $X=205890 $Y=176560
X2494 VSS VDD 339 364 339 269 ICV_41 $T=65320 165920 0 0 $X=65130 $Y=165680
X2495 VSS VDD 477 462 357 463 ICV_41 $T=87400 214880 1 0 $X=87210 $Y=211920
X2496 VSS VDD 624 624 690 685 ICV_41 $T=136620 182240 1 0 $X=136430 $Y=179280
X2497 VSS VDD 618 804 337 444 ICV_41 $T=160080 171360 0 0 $X=159890 $Y=171120
X2498 VSS VDD 894 894 769 882 ICV_41 $T=172500 149600 1 0 $X=172310 $Y=146640
X2499 VSS VDD 913 893 892 861 ICV_41 $T=175720 122400 0 0 $X=175530 $Y=122160
X2500 VSS VDD 1008 1008 784 999 ICV_41 $T=203320 62560 1 0 $X=203130 $Y=59600
X2501 VSS VDD 997 661 727 997 ICV_41 $T=206080 144160 1 0 $X=205890 $Y=141200
X2502 VSS VDD ICV_42 $T=6900 176800 1 0 $X=6710 $Y=173840
X2503 VSS VDD ICV_42 $T=6900 225760 0 0 $X=6710 $Y=225520
X2504 VSS VDD ICV_42 $T=18400 116960 0 0 $X=18210 $Y=116720
X2505 VSS VDD ICV_42 $T=20240 13600 1 0 $X=20050 $Y=10640
X2506 VSS VDD ICV_42 $T=20240 122400 1 0 $X=20050 $Y=119440
X2507 VSS VDD ICV_42 $T=20240 144160 1 0 $X=20050 $Y=141200
X2508 VSS VDD ICV_42 $T=24380 78880 1 0 $X=24190 $Y=75920
X2509 VSS VDD ICV_42 $T=33120 187680 1 0 $X=32930 $Y=184720
X2510 VSS VDD ICV_42 $T=34040 40800 0 0 $X=33850 $Y=40560
X2511 VSS VDD ICV_42 $T=37720 160480 0 0 $X=37530 $Y=160240
X2512 VSS VDD ICV_42 $T=48300 116960 1 0 $X=48110 $Y=114000
X2513 VSS VDD ICV_42 $T=50600 187680 1 0 $X=50410 $Y=184720
X2514 VSS VDD ICV_42 $T=64860 198560 1 0 $X=64670 $Y=195600
X2515 VSS VDD ICV_42 $T=73600 84320 0 0 $X=73410 $Y=84080
X2516 VSS VDD ICV_42 $T=77280 225760 0 0 $X=77090 $Y=225520
X2517 VSS VDD ICV_42 $T=80500 100640 1 0 $X=80310 $Y=97680
X2518 VSS VDD ICV_42 $T=85100 171360 1 0 $X=84910 $Y=168400
X2519 VSS VDD ICV_42 $T=85560 35360 1 0 $X=85370 $Y=32400
X2520 VSS VDD ICV_42 $T=89240 40800 1 0 $X=89050 $Y=37840
X2521 VSS VDD ICV_42 $T=104420 165920 1 0 $X=104230 $Y=162960
X2522 VSS VDD ICV_42 $T=118220 51680 0 0 $X=118030 $Y=51440
X2523 VSS VDD ICV_42 $T=120060 13600 1 0 $X=119870 $Y=10640
X2524 VSS VDD ICV_42 $T=120520 171360 1 0 $X=120330 $Y=168400
X2525 VSS VDD ICV_42 $T=121900 116960 0 0 $X=121710 $Y=116720
X2526 VSS VDD ICV_42 $T=130180 171360 0 0 $X=129990 $Y=171120
X2527 VSS VDD ICV_42 $T=137080 214880 1 0 $X=136890 $Y=211920
X2528 VSS VDD ICV_42 $T=141680 62560 1 0 $X=141490 $Y=59600
X2529 VSS VDD ICV_42 $T=145820 24480 1 0 $X=145630 $Y=21520
X2530 VSS VDD ICV_42 $T=145820 193120 1 0 $X=145630 $Y=190160
X2531 VSS VDD ICV_42 $T=160540 24480 1 0 $X=160350 $Y=21520
X2532 VSS VDD ICV_42 $T=160540 165920 1 0 $X=160350 $Y=162960
X2533 VSS VDD ICV_42 $T=160540 214880 1 0 $X=160350 $Y=211920
X2534 VSS VDD ICV_42 $T=162380 160480 0 0 $X=162190 $Y=160240
X2535 VSS VDD ICV_42 $T=167900 111520 1 0 $X=167710 $Y=108560
X2536 VSS VDD ICV_42 $T=174340 106080 0 0 $X=174150 $Y=105840
X2537 VSS VDD ICV_42 $T=177100 225760 0 0 $X=176910 $Y=225520
X2538 VSS VDD ICV_42 $T=178480 198560 0 0 $X=178290 $Y=198320
X2539 VSS VDD ICV_42 $T=180320 68000 0 0 $X=180130 $Y=67760
X2540 VSS VDD ICV_42 $T=188600 73440 1 0 $X=188410 $Y=70480
X2541 VSS VDD ICV_42 $T=205620 225760 0 0 $X=205430 $Y=225520
X2542 VSS VDD 20 94 270 ICV_43 $T=44620 133280 0 0 $X=44430 $Y=133040
X2543 VSS VDD 331 316 271 ICV_43 $T=54740 144160 0 0 $X=54550 $Y=143920
X2544 VSS VDD 362 43 387 ICV_43 $T=69000 68000 1 0 $X=68810 $Y=65040
X2545 VSS VDD 458 443 448 ICV_43 $T=82800 51680 0 0 $X=82610 $Y=51440
X2546 VSS VDD 425 331 418 ICV_43 $T=83260 149600 0 0 $X=83070 $Y=149360
X2547 VSS VDD 530 515 393 ICV_43 $T=97520 111520 1 0 $X=97330 $Y=108560
X2548 VSS VDD 551 527 542 ICV_43 $T=100740 68000 0 0 $X=100550 $Y=67760
X2549 VSS VDD 456 20 567 ICV_43 $T=104420 95200 0 0 $X=104230 $Y=94960
X2550 VSS VDD 586 516 516 ICV_43 $T=111320 13600 0 0 $X=111130 $Y=13360
X2551 VSS VDD 522 628 519 ICV_43 $T=118680 46240 1 0 $X=118490 $Y=43280
X2552 VSS VDD 629 509 650 ICV_43 $T=125580 84320 0 0 $X=125390 $Y=84080
X2553 VSS VDD 730 632 623 ICV_43 $T=133860 40800 0 0 $X=133670 $Y=40560
X2554 VSS VDD 736 716 726 ICV_43 $T=135240 95200 0 0 $X=135050 $Y=94960
X2555 VSS VDD 693 757 776 ICV_43 $T=147200 133280 1 0 $X=147010 $Y=130320
X2556 VSS VDD 755 766 766 ICV_43 $T=153640 133280 1 0 $X=153450 $Y=130320
X2557 VSS VDD 770 770 798 ICV_43 $T=153640 204000 1 0 $X=153450 $Y=201040
X2558 VSS VDD 876 596 861 ICV_43 $T=165600 116960 0 0 $X=165410 $Y=116720
X2559 VSS VDD 827 698 856 ICV_43 $T=166980 111520 0 0 $X=166790 $Y=111280
X2560 VSS VDD 885 815 875 ICV_43 $T=167440 51680 0 0 $X=167250 $Y=51440
X2561 VSS VDD 596 745 551 ICV_43 $T=167440 68000 0 0 $X=167250 $Y=67760
X2562 VSS VDD 547 905 896 ICV_43 $T=179400 182240 1 0 $X=179210 $Y=179280
X2563 VSS VDD 784 749 912 ICV_43 $T=181240 51680 1 0 $X=181050 $Y=48720
X2564 VSS VDD 946 914 914 ICV_43 $T=189520 182240 1 0 $X=189330 $Y=179280
X2565 VSS VDD 701 670 650 ICV_43 $T=193200 46240 1 0 $X=193010 $Y=43280
X2566 VSS VDD 776 928 973 ICV_43 $T=193200 127840 0 0 $X=193010 $Y=127600
X2567 VSS VDD 990 968 980 ICV_43 $T=193660 214880 0 0 $X=193470 $Y=214640
X2568 VSS VDD 960 SCAN_IN<2> SCAN_IN<3> ICV_43 $T=195500 193120 0 0 $X=195310 $Y=192880
X2569 VSS VDD 988 998 1031 ICV_43 $T=205620 149600 0 0 $X=205430 $Y=149360
X2570 VSS VDD 139 19 ICV_44 $T=20240 24480 1 0 $X=20050 $Y=21520
X2571 VSS VDD 174 118 ICV_44 $T=24840 160480 0 0 $X=24650 $Y=160240
X2572 VSS VDD 148 173 ICV_44 $T=25300 155040 0 0 $X=25110 $Y=154800
X2573 VSS VDD 489 502 ICV_44 $T=90160 46240 0 0 $X=89970 $Y=46000
X2574 VSS VDD 413 666 ICV_44 $T=120060 106080 0 0 $X=119870 $Y=105840
X2575 VSS VDD 684 608 ICV_44 $T=126500 35360 0 0 $X=126310 $Y=35120
X2576 VSS VDD 777 787 ICV_44 $T=146280 155040 0 0 $X=146090 $Y=154800
X2577 VSS VDD 660 16 ICV_44 $T=146280 209440 0 0 $X=146090 $Y=209200
X2578 VSS VDD 730 776 ICV_44 $T=155020 106080 0 0 $X=154830 $Y=105840
X2579 VSS VDD 818 821 ICV_44 $T=157780 13600 0 0 $X=157590 $Y=13360
X2580 VSS VDD 853 865 ICV_44 $T=163300 13600 0 0 $X=163110 $Y=13360
X2581 VSS VDD 1020 1028 ICV_44 $T=202860 24480 1 0 $X=202670 $Y=21520
X2582 VSS VDD 1014 1033 ICV_44 $T=204240 204000 0 0 $X=204050 $Y=203760
X2583 VSS VDD 996 995 ICV_44 $T=205620 84320 1 0 $X=205430 $Y=81360
X2584 VSS VDD 102 90 104 VDD 161 VSS sky130_fd_sc_hd__o21ai_4 $T=21160 176800 1 0 $X=20970 $Y=173840
X2585 VSS VDD 119 193 198 VDD 192 VSS sky130_fd_sc_hd__o21ai_4 $T=34040 73440 1 0 $X=33850 $Y=70480
X2586 VSS VDD 201 165 199 VDD 236 VSS sky130_fd_sc_hd__o21ai_4 $T=34960 89760 0 0 $X=34770 $Y=89520
X2587 VSS VDD 330 119 323 VDD 354 VSS sky130_fd_sc_hd__o21ai_4 $T=58420 73440 1 0 $X=58230 $Y=70480
X2588 VSS VDD 348 356 316 VDD 335 VSS sky130_fd_sc_hd__o21ai_4 $T=63480 155040 1 0 $X=63290 $Y=152080
X2589 VSS VDD 345 CLK_OUT 281 VDD 384 VSS sky130_fd_sc_hd__o21ai_4 $T=65780 100640 1 0 $X=65590 $Y=97680
X2590 VSS VDD 393 125 405 VDD 434 VSS sky130_fd_sc_hd__o21ai_4 $T=74520 78880 0 0 $X=74330 $Y=78640
X2591 VSS VDD 414 403 408 VDD 244 VSS sky130_fd_sc_hd__o21ai_4 $T=77280 176800 1 0 $X=77090 $Y=173840
X2592 VSS VDD 428 406 436 VDD 195 VSS sky130_fd_sc_hd__o21ai_4 $T=78200 133280 0 0 $X=78010 $Y=133040
X2593 VSS VDD 378 410 444 VDD 403 VSS sky130_fd_sc_hd__o21ai_4 $T=78660 171360 0 0 $X=78470 $Y=171120
X2594 VSS VDD 565 570 577 VDD 622 VSS sky130_fd_sc_hd__o21ai_4 $T=111780 57120 1 0 $X=111590 $Y=54160
X2595 VSS VDD 658 652 648 VDD 599 VSS sky130_fd_sc_hd__o21ai_4 $T=123280 100640 0 0 $X=123090 $Y=100400
X2596 VSS VDD 717 746 704 VDD 742 VSS sky130_fd_sc_hd__o21ai_4 $T=141220 116960 1 0 $X=141030 $Y=114000
X2597 VSS VDD 666 764 807 VDD 821 VSS sky130_fd_sc_hd__o21ai_4 $T=157320 19040 0 0 $X=157130 $Y=18800
X2598 VSS VDD 620 834 829 VDD 862 VSS sky130_fd_sc_hd__o21ai_4 $T=165600 187680 1 0 $X=165410 $Y=184720
X2599 VSS VDD 865 756 884 VDD 874 VSS sky130_fd_sc_hd__o21ai_4 $T=175260 35360 0 0 $X=175070 $Y=35120
X2600 VSS VDD 481 932 916 VDD 895 VSS sky130_fd_sc_hd__o21ai_4 $T=182160 171360 0 0 $X=181970 $Y=171120
X2601 VSS VDD 875 930 842 VDD 962 VSS sky130_fd_sc_hd__o21ai_4 $T=189520 35360 1 0 $X=189330 $Y=32400
X2602 VSS VDD 752 965 948 VDD 980 VSS sky130_fd_sc_hd__o21ai_4 $T=190900 204000 0 0 $X=190710 $Y=203760
X2603 VSS VDD 888 932 950 VDD 986 VSS sky130_fd_sc_hd__o21ai_4 $T=192280 89760 0 0 $X=192090 $Y=89520
X2604 VSS VDD 967 965 961 VDD 1007 VSS sky130_fd_sc_hd__o21ai_4 $T=196420 193120 1 0 $X=196230 $Y=190160
X2605 VSS VDD 957 1011 1010 VDD 907 VSS sky130_fd_sc_hd__o21ai_4 $T=205160 220320 1 0 $X=204970 $Y=217360
X2606 VSS VDD ICV_45 $T=23000 220320 0 0 $X=22810 $Y=220080
X2607 VSS VDD ICV_45 $T=40940 193120 1 0 $X=40750 $Y=190160
X2608 VSS VDD ICV_45 $T=52440 165920 1 0 $X=52250 $Y=162960
X2609 VSS VDD ICV_45 $T=104420 62560 1 0 $X=104230 $Y=59600
X2610 VSS VDD ICV_45 $T=111780 46240 1 0 $X=111590 $Y=43280
X2611 VSS VDD ICV_45 $T=134780 24480 1 0 $X=134590 $Y=21520
X2612 VSS VDD ICV_45 $T=137540 73440 1 0 $X=137350 $Y=70480
X2613 VSS VDD ICV_45 $T=137540 138720 1 0 $X=137350 $Y=135760
X2614 VSS VDD ICV_45 $T=163300 19040 0 0 $X=163110 $Y=18800
X2615 VSS VDD ICV_45 $T=164220 106080 1 0 $X=164030 $Y=103120
X2616 VSS VDD ICV_45 $T=191360 84320 0 0 $X=191170 $Y=84080
X2617 VSS VDD ICV_45 $T=196420 62560 1 0 $X=196230 $Y=59600
X2618 VSS VDD ICV_45 $T=205160 165920 1 0 $X=204970 $Y=162960
X2619 VSS VDD 136 93 ICV_46 $T=20240 127840 1 0 $X=20050 $Y=124880
X2620 VSS VDD SCAN_IN<21> 95 ICV_46 $T=34040 133280 0 0 $X=33850 $Y=133040
X2621 VSS VDD 383 391 ICV_46 $T=80040 29920 0 0 $X=79850 $Y=29680
X2622 VSS VDD 472 478 ICV_46 $T=86480 127840 1 0 $X=86290 $Y=124880
X2623 VSS VDD 572 529 ICV_46 $T=104880 62560 0 0 $X=104690 $Y=62320
X2624 VSS VDD 796 796 ICV_46 $T=153640 29920 1 0 $X=153450 $Y=26960
X2625 VSS VDD 899 900 ICV_46 $T=170660 127840 1 0 $X=170470 $Y=124880
X2626 VSS VDD 950 888 ICV_46 $T=186300 89760 0 0 $X=186110 $Y=89520
X2627 VSS VDD 1029 158 ICV_46 $T=205160 111520 1 0 $X=204970 $Y=108560
X2628 VSS VDD 95 114 114 ICV_47 $T=20700 149600 0 0 $X=20510 $Y=149360
X2629 VSS VDD 307 261 261 ICV_47 $T=46000 46240 0 0 $X=45810 $Y=46000
X2630 VSS VDD 294 250 287 ICV_47 $T=47840 35360 0 0 $X=47650 $Y=35120
X2631 VSS VDD 255 285 285 ICV_47 $T=49220 95200 0 0 $X=49030 $Y=94960
X2632 VSS VDD 361 383 383 ICV_47 $T=69460 35360 0 0 $X=69270 $Y=35120
X2633 VSS VDD 449 SCAN_IN<20> 498 ICV_47 $T=92460 116960 1 0 $X=92270 $Y=114000
X2634 VSS VDD 604 510 510 ICV_47 $T=105800 51680 0 0 $X=105610 $Y=51440
X2635 VSS VDD 775 674 608 ICV_47 $T=146280 29920 0 0 $X=146090 $Y=29680
X2636 VSS VDD 1044 984 1016 ICV_47 $T=204700 176800 1 0 $X=204510 $Y=173840
X2637 VSS VDD 145 141 65 VDD 123 VSS sky130_fd_sc_hd__o21a_4 $T=21620 204000 0 0 $X=21430 $Y=203760
X2638 VSS VDD 140 120 159 VDD 165 VSS sky130_fd_sc_hd__o21a_4 $T=27140 106080 1 0 $X=26950 $Y=103120
X2639 VSS VDD 143 87 132 VDD 144 VSS sky130_fd_sc_hd__o21a_4 $T=27600 187680 1 0 $X=27410 $Y=184720
X2640 VSS VDD 170 147 139 VDD 169 VSS sky130_fd_sc_hd__o21a_4 $T=28060 19040 1 0 $X=27870 $Y=16080
X2641 VSS VDD 182 168 157 VDD 185 VSS sky130_fd_sc_hd__o21a_4 $T=31740 51680 1 0 $X=31550 $Y=48720
X2642 VSS VDD 196 200 219 VDD 174 VSS sky130_fd_sc_hd__o21a_4 $T=34960 160480 1 0 $X=34770 $Y=157520
X2643 VSS VDD 176 SCAN_IN<21> 102 VDD 206 VSS sky130_fd_sc_hd__o21a_4 $T=34960 182240 1 0 $X=34770 $Y=179280
X2644 VSS VDD 242 255 217 VDD 211 VSS sky130_fd_sc_hd__o21a_4 $T=43700 95200 0 0 $X=43510 $Y=94960
X2645 VSS VDD 272 282 301 VDD 146 VSS sky130_fd_sc_hd__o21a_4 $T=50140 209440 0 0 $X=49950 $Y=209200
X2646 VSS VDD 145 305 280 VDD 291 VSS sky130_fd_sc_hd__o21a_4 $T=50140 220320 1 0 $X=49950 $Y=217360
X2647 VSS VDD 286 310 338 VDD 340 VSS sky130_fd_sc_hd__o21a_4 $T=61180 182240 1 0 $X=60990 $Y=179280
X2648 VSS VDD 346 321 248 VDD 293 VSS sky130_fd_sc_hd__o21a_4 $T=63020 171360 0 0 $X=62830 $Y=171120
X2649 VSS VDD 238 386 397 VDD 312 VSS sky130_fd_sc_hd__o21a_4 $T=71760 24480 0 0 $X=71570 $Y=24240
X2650 VSS VDD 213 300 426 VDD 419 VSS sky130_fd_sc_hd__o21a_4 $T=77280 193120 1 0 $X=77090 $Y=190160
X2651 VSS VDD 92 415 301 VDD 374 VSS sky130_fd_sc_hd__o21a_4 $T=77280 214880 1 0 $X=77090 $Y=211920
X2652 VSS VDD 448 471 248 VDD 468 VSS sky130_fd_sc_hd__o21a_4 $T=88320 149600 1 0 $X=88130 $Y=146640
X2653 VSS VDD 433 481 499 VDD 451 VSS sky130_fd_sc_hd__o21a_4 $T=93840 176800 1 0 $X=93650 $Y=173840
X2654 VSS VDD 501 489 502 VDD 452 VSS sky130_fd_sc_hd__o21a_4 $T=94760 51680 1 0 $X=94570 $Y=48720
X2655 VSS VDD 531 SCAN_IN<19> 247 VDD 518 VSS sky130_fd_sc_hd__o21a_4 $T=98900 122400 0 0 $X=98710 $Y=122160
X2656 VSS VDD 357 492 583 VDD 544 VSS sky130_fd_sc_hd__o21a_4 $T=104420 220320 0 0 $X=104230 $Y=220080
X2657 VSS VDD 472 494 517 VDD 555 VSS sky130_fd_sc_hd__o21a_4 $T=105340 133280 1 0 $X=105150 $Y=130320
X2658 VSS VDD 566 SCAN_IN<21> 565 VDD 578 VSS sky130_fd_sc_hd__o21a_4 $T=108560 89760 1 0 $X=108370 $Y=86800
X2659 VSS VDD 92 579 301 VDD 595 VSS sky130_fd_sc_hd__o21a_4 $T=111320 214880 1 0 $X=111130 $Y=211920
X2660 VSS VDD 608 609 591 VDD 571 VSS sky130_fd_sc_hd__o21a_4 $T=115920 35360 1 0 $X=115730 $Y=32400
X2661 VSS VDD 638 529 607 VDD 548 VSS sky130_fd_sc_hd__o21a_4 $T=119140 62560 0 0 $X=118950 $Y=62320
X2662 VSS VDD 550 641 646 VDD 515 VSS sky130_fd_sc_hd__o21a_4 $T=122820 198560 0 0 $X=122630 $Y=198320
X2663 VSS VDD 393 661 548 VDD 659 VSS sky130_fd_sc_hd__o21a_4 $T=123740 111520 0 0 $X=123550 $Y=111280
X2664 VSS VDD 649 707 695 VDD 687 VSS sky130_fd_sc_hd__o21a_4 $T=133400 51680 1 0 $X=133210 $Y=48720
X2665 VSS VDD 393 698 548 VDD 689 VSS sky130_fd_sc_hd__o21a_4 $T=133400 84320 1 0 $X=133210 $Y=81360
X2666 VSS VDD 691 665 682 VDD 715 VSS sky130_fd_sc_hd__o21a_4 $T=135700 187680 0 0 $X=135510 $Y=187440
X2667 VSS VDD 731 453 745 VDD 684 VSS sky130_fd_sc_hd__o21a_4 $T=137540 68000 1 0 $X=137350 $Y=65040
X2668 VSS VDD 722 721 733 VDD 737 VSS sky130_fd_sc_hd__o21a_4 $T=139380 127840 1 0 $X=139190 $Y=124880
X2669 VSS VDD 509 759 769 VDD 718 VSS sky130_fd_sc_hd__o21a_4 $T=143060 149600 1 0 $X=142870 $Y=146640
X2670 VSS VDD 786 633 537 VDD 682 VSS sky130_fd_sc_hd__o21a_4 $T=148580 198560 1 0 $X=148390 $Y=195600
X2671 VSS VDD 608 780 775 VDD 781 VSS sky130_fd_sc_hd__o21a_4 $T=150880 35360 1 0 $X=150690 $Y=32400
X2672 VSS VDD 783 791 785 VDD 800 VSS sky130_fd_sc_hd__o21a_4 $T=156400 149600 0 0 $X=156210 $Y=149360
X2673 VSS VDD 551 592 745 VDD 808 VSS sky130_fd_sc_hd__o21a_4 $T=157780 116960 0 0 $X=157590 $Y=116720
X2674 VSS VDD 513 788 815 VDD 443 VSS sky130_fd_sc_hd__o21a_4 $T=161000 46240 0 0 $X=160810 $Y=46000
X2675 VSS VDD 551 454 745 VDD 817 VSS sky130_fd_sc_hd__o21a_4 $T=161000 68000 0 0 $X=160810 $Y=67760
X2676 VSS VDD 840 841 862 VDD 414 VSS sky130_fd_sc_hd__o21a_4 $T=164220 182240 0 0 $X=164030 $Y=182000
X2677 VSS VDD 885 888 921 VDD 503 VSS sky130_fd_sc_hd__o21a_4 $T=176180 84320 1 0 $X=175990 $Y=81360
X2678 VSS VDD 919 892 909 VDD 530 VSS sky130_fd_sc_hd__o21a_4 $T=178940 111520 0 0 $X=178750 $Y=111280
X2679 VSS VDD 1010 671 1014 VDD 992 VSS sky130_fd_sc_hd__o21a_4 $T=204240 214880 1 0 $X=204050 $Y=211920
X2680 VSS VDD 23 10 ICV_48 $T=7820 51680 1 0 $X=7630 $Y=48720
X2681 VSS VDD 16 52 ICV_48 $T=7820 204000 1 0 $X=7630 $Y=201040
X2682 VSS VDD 20 178 ICV_48 $T=34960 29920 0 0 $X=34770 $Y=29680
X2683 VSS VDD 199 239 ICV_48 $T=40020 78880 0 0 $X=39830 $Y=78640
X2684 VSS VDD 278 281 ICV_48 $T=49220 122400 1 0 $X=49030 $Y=119440
X2685 VSS VDD SCAN_IN<8> 263 ICV_48 $T=52900 149600 0 0 $X=52710 $Y=149360
X2686 VSS VDD 346 286 ICV_48 $T=62100 176800 1 0 $X=61910 $Y=173840
X2687 VSS VDD 295 358 ICV_48 $T=63020 133280 1 0 $X=62830 $Y=130320
X2688 VSS VDD CLK_OUT 345 ICV_48 $T=65780 95200 1 0 $X=65590 $Y=92240
X2689 VSS VDD 363 356 ICV_48 $T=69460 138720 0 0 $X=69270 $Y=138480
X2690 VSS VDD 379 391 ICV_48 $T=77280 46240 1 0 $X=77090 $Y=43280
X2691 VSS VDD 231 436 ICV_48 $T=78200 133280 1 0 $X=78010 $Y=130320
X2692 VSS VDD 240 460 ICV_48 $T=84640 204000 0 0 $X=84450 $Y=203760
X2693 VSS VDD 20 416 ICV_48 $T=92920 111520 1 0 $X=92730 $Y=108560
X2694 VSS VDD 492 583 ICV_48 $T=110860 220320 0 0 $X=110670 $Y=220080
X2695 VSS VDD 624 485 ICV_48 $T=118220 133280 1 0 $X=118030 $Y=130320
X2696 VSS VDD 625 458 ICV_48 $T=118220 160480 1 0 $X=118030 $Y=157520
X2697 VSS VDD SCAN_IN<11> 661 ICV_48 $T=132480 111520 0 0 $X=132290 $Y=111280
X2698 VSS VDD 690 624 ICV_48 $T=137080 176800 0 0 $X=136890 $Y=176560
X2699 VSS VDD 728 738 ICV_48 $T=137080 198560 0 0 $X=136890 $Y=198320
X2700 VSS VDD 710 742 ICV_48 $T=138920 95200 1 0 $X=138730 $Y=92240
X2701 VSS VDD 673 673 ICV_48 $T=138920 165920 0 0 $X=138730 $Y=165680
X2702 VSS VDD 704 746 ICV_48 $T=142140 111520 1 0 $X=141950 $Y=108560
X2703 VSS VDD 744 773 ICV_48 $T=146280 40800 1 0 $X=146090 $Y=37840
X2704 VSS VDD 760 760 ICV_48 $T=147660 160480 1 0 $X=147470 $Y=157520
X2705 VSS VDD 817 824 ICV_48 $T=160080 62560 0 0 $X=159890 $Y=62320
X2706 VSS VDD 738 798 ICV_48 $T=160540 187680 0 0 $X=160350 $Y=187440
X2707 VSS VDD 810 802 ICV_48 $T=162840 51680 0 0 $X=162650 $Y=51440
X2708 VSS VDD 810 790 ICV_48 $T=168820 57120 0 0 $X=168630 $Y=56880
X2709 VSS VDD 892 900 ICV_48 $T=176180 122400 1 0 $X=175990 $Y=119440
X2710 VSS VDD 885 875 ICV_48 $T=176640 51680 1 0 $X=176450 $Y=48720
X2711 VSS VDD SCAN_IN<7> 887 ICV_48 $T=180320 13600 0 0 $X=180130 $Y=13360
X2712 VSS VDD 924 931 ICV_48 $T=180320 165920 0 0 $X=180130 $Y=165680
X2713 VSS VDD 769 940 ICV_48 $T=183080 144160 1 0 $X=182890 $Y=141200
X2714 VSS VDD 995 914 ICV_48 $T=200560 100640 1 0 $X=200370 $Y=97680
X2715 VSS VDD 727 1005 ICV_48 $T=203780 171360 1 0 $X=203590 $Y=168400
X2716 VSS VDD 33 79 ICV_49 $T=12420 204000 1 0 $X=12230 $Y=201040
X2717 VSS VDD 224 262 ICV_49 $T=49220 46240 1 0 $X=49030 $Y=43280
X2718 VSS VDD 458 503 ICV_49 $T=92920 89760 1 0 $X=92730 $Y=86800
X2719 VSS VDD 550 590 ICV_49 $T=112240 176800 0 0 $X=112050 $Y=176560
X2720 VSS VDD 787 771 ICV_49 $T=166060 78880 0 0 $X=165870 $Y=78640
X2721 VSS VDD 866 825 ICV_49 $T=167900 73440 0 0 $X=167710 $Y=73200
X2722 VSS VDD 889 907 ICV_49 $T=174800 209440 1 0 $X=174610 $Y=206480
X2723 VSS VDD 752 965 ICV_49 $T=190900 204000 1 0 $X=190710 $Y=201040
X2724 VSS VDD 20 844 ICV_49 $T=203780 78880 1 0 $X=203590 $Y=75920
X2725 VSS VDD 20 53 ICV_50 $T=7820 29920 1 0 $X=7630 $Y=26960
X2726 VSS VDD 164 181 ICV_50 $T=34960 68000 0 0 $X=34770 $Y=67760
X2727 VSS VDD 356 438 ICV_50 $T=79580 116960 1 0 $X=79390 $Y=114000
X2728 VSS VDD 410 444 ICV_50 $T=85560 171360 0 0 $X=85370 $Y=171120
X2729 VSS VDD 190 546 ICV_50 $T=112700 187680 1 0 $X=112510 $Y=184720
X2730 VSS VDD 621 627 ICV_50 $T=116380 209440 1 0 $X=116190 $Y=206480
X2731 VSS VDD 714 735 ICV_50 $T=136620 29920 0 0 $X=136430 $Y=29680
X2732 VSS VDD 759 790 ICV_50 $T=152260 144160 0 0 $X=152070 $Y=143920
X2733 VSS VDD 904 666 ICV_50 $T=184460 57120 0 0 $X=184270 $Y=56880
X2734 VSS VDD 823 SCAN_IN<3> ICV_50 $T=186760 204000 0 0 $X=186570 $Y=203760
X2735 VSS VDD 992 980 ICV_50 $T=197800 204000 0 0 $X=197610 $Y=203760
X2736 VSS VDD 701 985 ICV_50 $T=201020 68000 1 0 $X=200830 $Y=65040
X2737 VSS VDD 940 1003 ICV_50 $T=203320 106080 0 0 $X=203130 $Y=105840
X2738 VSS VDD 44 ICV_51 $T=6900 78880 1 0 $X=6710 $Y=75920
X2739 VSS VDD 55 ICV_51 $T=6900 84320 1 0 $X=6710 $Y=81360
X2740 VSS VDD 81 ICV_51 $T=17480 57120 0 0 $X=17290 $Y=56880
X2741 VSS VDD 500 ICV_51 $T=92000 204000 0 0 $X=91810 $Y=203760
X2742 VSS VDD 609 ICV_51 $T=111320 35360 1 0 $X=111130 $Y=32400
X2743 VSS VDD 637 ICV_51 $T=117300 40800 1 0 $X=117110 $Y=37840
X2744 VSS VDD 646 ICV_51 $T=118220 198560 0 0 $X=118030 $Y=198320
X2745 VSS VDD 290 ICV_51 $T=118220 209440 0 0 $X=118030 $Y=209200
X2746 VSS VDD 619 ICV_51 $T=121900 182240 0 0 $X=121710 $Y=182000
X2747 VSS VDD 670 ICV_51 $T=123280 68000 0 0 $X=123090 $Y=67760
X2748 VSS VDD 974 ICV_51 $T=191360 13600 1 0 $X=191170 $Y=10640
X2749 VSS VDD 1019 ICV_51 $T=202400 100640 0 0 $X=202210 $Y=100400
X2750 VSS VDD 960 ICV_51 $T=202400 198560 0 0 $X=202210 $Y=198320
X2751 VSS 353 ICV_52 $T=61640 176800 0 0 $X=61450 $Y=176560
X2752 VSS 424 ICV_52 $T=75900 182240 1 0 $X=75710 $Y=179280
X2753 VSS 448 ICV_52 $T=89700 84320 0 0 $X=89510 $Y=84080
X2754 VSS 481 ICV_52 $T=89700 193120 0 0 $X=89510 $Y=192880
X2755 VSS 245 ICV_52 $T=89700 204000 0 0 $X=89510 $Y=203760
X2756 VSS 462 ICV_52 $T=89700 209440 0 0 $X=89510 $Y=209200
X2757 VSS 598 ICV_52 $T=117760 100640 0 0 $X=117570 $Y=100400
X2758 VSS SCAN_IN<16> ICV_52 $T=117760 106080 0 0 $X=117570 $Y=105840
X2759 VSS 688 ICV_52 $T=132020 68000 1 0 $X=131830 $Y=65040
X2760 VSS 618 ICV_52 $T=132020 160480 1 0 $X=131830 $Y=157520
X2761 VSS 731 ICV_52 $T=145820 68000 0 0 $X=145630 $Y=67760
X2762 VSS 899 ICV_52 $T=173880 133280 0 0 $X=173690 $Y=133040
X2763 VSS 901 ICV_52 $T=188140 225760 1 0 $X=187950 $Y=222800
X2764 VSS 980 ICV_52 $T=201940 204000 0 0 $X=201750 $Y=203760
X2765 VSS VDD ICV_53 $T=19780 29920 1 0 $X=19590 $Y=26960
X2766 VSS VDD ICV_53 $T=19780 106080 1 0 $X=19590 $Y=103120
X2767 VSS VDD ICV_53 $T=19780 149600 1 0 $X=19590 $Y=146640
X2768 VSS VDD ICV_53 $T=33580 171360 0 0 $X=33390 $Y=171120
X2769 VSS VDD ICV_53 $T=34040 13600 1 0 $X=33850 $Y=10640
X2770 VSS VDD ICV_53 $T=47840 193120 1 0 $X=47650 $Y=190160
X2771 VSS VDD ICV_53 $T=61640 57120 0 0 $X=61450 $Y=56880
X2772 VSS VDD ICV_53 $T=75900 220320 1 0 $X=75710 $Y=217360
X2773 VSS VDD ICV_53 $T=89700 51680 0 0 $X=89510 $Y=51440
X2774 VSS VDD ICV_53 $T=89700 149600 0 0 $X=89510 $Y=149360
X2775 VSS VDD ICV_53 $T=89700 171360 0 0 $X=89510 $Y=171120
X2776 VSS VDD ICV_53 $T=103960 24480 1 0 $X=103770 $Y=21520
X2777 VSS VDD ICV_53 $T=103960 78880 1 0 $X=103770 $Y=75920
X2778 VSS VDD ICV_53 $T=103960 106080 1 0 $X=103770 $Y=103120
X2779 VSS VDD ICV_53 $T=103960 111520 1 0 $X=103770 $Y=108560
X2780 VSS VDD ICV_53 $T=103960 116960 1 0 $X=103770 $Y=114000
X2781 VSS VDD ICV_53 $T=103960 144160 1 0 $X=103770 $Y=141200
X2782 VSS VDD ICV_53 $T=117760 89760 0 0 $X=117570 $Y=89520
X2783 VSS VDD ICV_53 $T=132020 133280 1 0 $X=131830 $Y=130320
X2784 VSS VDD ICV_53 $T=132020 149600 1 0 $X=131830 $Y=146640
X2785 VSS VDD ICV_53 $T=132020 165920 1 0 $X=131830 $Y=162960
X2786 VSS VDD ICV_53 $T=145820 100640 0 0 $X=145630 $Y=100400
X2787 VSS VDD ICV_53 $T=145820 149600 0 0 $X=145630 $Y=149360
X2788 VSS VDD ICV_53 $T=173880 89760 0 0 $X=173690 $Y=89520
X2789 VSS VDD ICV_53 $T=173880 160480 0 0 $X=173690 $Y=160240
X2790 VSS VDD ICV_53 $T=173880 171360 0 0 $X=173690 $Y=171120
X2791 VSS VDD ICV_53 $T=188140 46240 1 0 $X=187950 $Y=43280
X2792 VSS VDD ICV_53 $T=188140 84320 1 0 $X=187950 $Y=81360
X2793 VSS VDD ICV_53 $T=188140 116960 1 0 $X=187950 $Y=114000
X2794 VSS VDD ICV_53 $T=188140 122400 1 0 $X=187950 $Y=119440
X2795 VSS VDD ICV_53 $T=188140 144160 1 0 $X=187950 $Y=141200
X2796 VSS VDD ICV_53 $T=190900 225760 0 0 $X=190710 $Y=225520
X2797 VSS VDD ICV_53 $T=201940 24480 0 0 $X=201750 $Y=24240
X2798 VSS VDD ICV_53 $T=201940 29920 0 0 $X=201750 $Y=29680
X2799 VSS VDD ICV_53 $T=201940 176800 0 0 $X=201750 $Y=176560
X2800 VSS VDD ICV_53 $T=201940 182240 0 0 $X=201750 $Y=182000
X2801 VSS VDD ICV_54 $T=33580 24480 0 0 $X=33390 $Y=24240
X2802 VSS VDD ICV_54 $T=47840 19040 1 0 $X=47650 $Y=16080
X2803 VSS VDD ICV_54 $T=47840 57120 1 0 $X=47650 $Y=54160
X2804 VSS VDD ICV_54 $T=47840 62560 1 0 $X=47650 $Y=59600
X2805 VSS VDD ICV_54 $T=47840 100640 1 0 $X=47650 $Y=97680
X2806 VSS VDD ICV_54 $T=89700 89760 0 0 $X=89510 $Y=89520
X2807 VSS VDD ICV_54 $T=103960 95200 1 0 $X=103770 $Y=92240
X2808 VSS VDD ICV_54 $T=103960 122400 1 0 $X=103770 $Y=119440
X2809 VSS VDD ICV_54 $T=132020 209440 1 0 $X=131830 $Y=206480
X2810 VSS VDD ICV_54 $T=132020 214880 1 0 $X=131830 $Y=211920
X2811 VSS VDD ICV_54 $T=132020 225760 1 0 $X=131830 $Y=222800
X2812 VSS VDD ICV_54 $T=145820 13600 0 0 $X=145630 $Y=13360
X2813 VSS VDD ICV_54 $T=160080 149600 1 0 $X=159890 $Y=146640
X2814 VSS VDD ICV_54 $T=160080 182240 1 0 $X=159890 $Y=179280
X2815 VSS VDD ICV_54 $T=173880 122400 0 0 $X=173690 $Y=122160
X2816 VSS VDD ICV_54 $T=173880 127840 0 0 $X=173690 $Y=127600
X2817 VSS VDD ICV_54 $T=173880 187680 0 0 $X=173690 $Y=187440
X2818 VSS VDD ICV_54 $T=201940 89760 0 0 $X=201750 $Y=89520
X2819 VSS VDD ICV_54 $T=201940 165920 0 0 $X=201750 $Y=165680
X2820 VSS VDD ICV_55 $T=19780 35360 1 0 $X=19590 $Y=32400
X2821 VSS VDD ICV_55 $T=33580 187680 0 0 $X=33390 $Y=187440
X2822 VSS VDD ICV_55 $T=47840 84320 1 0 $X=47650 $Y=81360
X2823 VSS VDD ICV_55 $T=47840 95200 1 0 $X=47650 $Y=92240
X2824 VSS VDD ICV_55 $T=61640 187680 0 0 $X=61450 $Y=187440
X2825 VSS VDD ICV_55 $T=75900 68000 1 0 $X=75710 $Y=65040
X2826 VSS VDD ICV_55 $T=89700 40800 0 0 $X=89510 $Y=40560
X2827 VSS VDD ICV_55 $T=103960 35360 1 0 $X=103770 $Y=32400
X2828 VSS VDD ICV_55 $T=105340 225760 0 0 $X=105150 $Y=225520
X2829 VSS VDD ICV_55 $T=132020 29920 1 0 $X=131830 $Y=26960
X2830 VSS VDD ICV_55 $T=132020 204000 1 0 $X=131830 $Y=201040
X2831 VSS VDD ICV_55 $T=201940 155040 0 0 $X=201750 $Y=154800
X2832 VSS VDD 116 70 ICV_56 $T=19780 19040 1 0 $X=19590 $Y=16080
X2833 VSS VDD 95 102 ICV_56 $T=33580 144160 0 0 $X=33390 $Y=143920
X2834 VSS VDD 187 118 ICV_56 $T=33580 165920 0 0 $X=33390 $Y=165680
X2835 VSS VDD 161 245 ICV_56 $T=47840 204000 1 0 $X=47650 $Y=201040
X2836 VSS VDD 225 290 ICV_56 $T=47840 214880 1 0 $X=47650 $Y=211920
X2837 VSS VDD 283 138 ICV_56 $T=47840 225760 1 0 $X=47650 $Y=222800
X2838 VSS VDD 327 315 ICV_56 $T=61640 144160 0 0 $X=61450 $Y=143920
X2839 VSS VDD 348 310 ICV_56 $T=61640 182240 0 0 $X=61450 $Y=182000
X2840 VSS VDD 390 147 ICV_56 $T=75900 19040 1 0 $X=75710 $Y=16080
X2841 VSS VDD 356 378 ICV_56 $T=75900 165920 1 0 $X=75710 $Y=162960
X2842 VSS VDD 420 301 ICV_56 $T=75900 225760 1 0 $X=75710 $Y=222800
X2843 VSS VDD 532 506 ICV_56 $T=103960 171360 1 0 $X=103770 $Y=168400
X2844 VSS VDD 672 632 ICV_56 $T=132020 95200 1 0 $X=131830 $Y=92240
X2845 VSS VDD 622 755 ICV_56 $T=145820 57120 0 0 $X=145630 $Y=56880
X2846 VSS VDD 578 766 ICV_56 $T=145820 62560 0 0 $X=145630 $Y=62320
X2847 VSS VDD 731 551 ICV_56 $T=145820 73440 0 0 $X=145630 $Y=73200
X2848 VSS VDD 767 736 ICV_56 $T=145820 89760 0 0 $X=145630 $Y=89520
X2849 VSS VDD 750 624 ICV_56 $T=145820 171360 0 0 $X=145630 $Y=171120
X2850 VSS VDD 618 568 ICV_56 $T=160080 176800 1 0 $X=159890 $Y=173840
X2851 VSS VDD 795 738 ICV_56 $T=160080 204000 1 0 $X=159890 $Y=201040
X2852 VSS VDD 882 791 ICV_56 $T=173880 155040 0 0 $X=173690 $Y=154800
X2853 VSS VDD 953 810 ICV_56 $T=188140 29920 1 0 $X=187950 $Y=26960
X2854 VSS VDD 911 771 ICV_56 $T=188140 51680 1 0 $X=187950 $Y=48720
X2855 VSS VDD 915 759 ICV_56 $T=188140 149600 1 0 $X=187950 $Y=146640
X2856 VSS VDD 998 661 ICV_56 $T=201940 149600 0 0 $X=201750 $Y=149360
X2857 VSS VDD 55 179 ICV_57 $T=33580 78880 0 0 $X=33390 $Y=78640
X2858 VSS VDD 345 421 ICV_57 $T=75900 95200 1 0 $X=75710 $Y=92240
X2859 VSS VDD 325 441 ICV_57 $T=89700 165920 0 0 $X=89510 $Y=165680
X2860 VSS VDD 615 605 ICV_57 $T=117760 122400 0 0 $X=117570 $Y=122160
X2861 VSS VDD 637 666 ICV_57 $T=132020 57120 1 0 $X=131830 $Y=54160
X2862 VSS VDD 878 887 ICV_57 $T=173880 13600 0 0 $X=173690 $Y=13360
X2863 VSS VDD 915 872 ICV_57 $T=173880 165920 0 0 $X=173690 $Y=165680
X2864 VSS VDD 972 977 ICV_57 $T=201940 116960 0 0 $X=201750 $Y=116720
X2865 VSS 173 196 ICV_58 $T=33580 160480 0 0 $X=33390 $Y=160240
X2866 VSS 251 361 ICV_58 $T=61640 29920 0 0 $X=61450 $Y=29680
X2867 VSS 128 350 ICV_58 $T=61640 40800 0 0 $X=61450 $Y=40560
X2868 VSS 276 26 ICV_58 $T=61640 78880 0 0 $X=61450 $Y=78640
X2869 VSS 58 491 ICV_58 $T=89700 198560 0 0 $X=89510 $Y=198320
X2870 VSS 442 492 ICV_58 $T=89700 220320 0 0 $X=89510 $Y=220080
X2871 VSS 535 543 ICV_58 $T=103960 198560 1 0 $X=103770 $Y=195600
X2872 VSS 549 507 ICV_58 $T=117760 149600 0 0 $X=117570 $Y=149360
X2873 VSS 395 645 ICV_58 $T=117760 182240 0 0 $X=117570 $Y=182000
X2874 VSS 696 646 ICV_58 $T=132020 198560 1 0 $X=131830 $Y=195600
X2875 VSS 16 20 ICV_58 $T=145820 214880 0 0 $X=145630 $Y=214640
X2876 VSS 697 724 ICV_58 $T=148120 13600 1 0 $X=147930 $Y=10640
X2877 VSS 892 909 ICV_58 $T=173880 111520 0 0 $X=173690 $Y=111280
X2878 VSS 784 955 ICV_58 $T=188140 62560 1 0 $X=187950 $Y=59600
X2879 VSS 1008 963 ICV_58 $T=201940 62560 0 0 $X=201750 $Y=62320
X2880 VSS VDD 172 179 ICV_59 $T=33580 84320 0 0 $X=33390 $Y=84080
X2881 VSS VDD 471 SCAN_IN<11> ICV_59 $T=89700 127840 0 0 $X=89510 $Y=127600
X2882 VSS VDD 708 708 ICV_59 $T=132020 220320 1 0 $X=131830 $Y=217360
X2883 VSS VDD 755 723 ICV_59 $T=145820 138720 0 0 $X=145630 $Y=138480
X2884 VSS VDD 829 841 ICV_59 $T=160080 187680 1 0 $X=159890 $Y=184720
X2885 VSS VDD 904 911 ICV_59 $T=173880 57120 0 0 $X=173690 $Y=56880
X2886 VSS VDD 847 17 ICV_59 $T=173880 73440 0 0 $X=173690 $Y=73200
X2887 VSS VDD 985 20 ICV_59 $T=201940 51680 0 0 $X=201750 $Y=51440
X2888 VSS VDD 43 55 112 ICV_60 $T=19780 78880 1 0 $X=19590 $Y=75920
X2889 VSS VDD 138 127 115 ICV_60 $T=33580 214880 0 0 $X=33390 $Y=214640
X2890 VSS VDD 162 202 183 ICV_60 $T=33580 220320 0 0 $X=33390 $Y=220080
X2891 VSS VDD 327 271 316 ICV_60 $T=61640 149600 0 0 $X=61450 $Y=149360
X2892 VSS VDD 289 330 379 ICV_60 $T=75900 57120 1 0 $X=75710 $Y=54160
X2893 VSS VDD 417 281 405 ICV_60 $T=75900 84320 1 0 $X=75710 $Y=81360
X2894 VSS VDD 535 547 500 ICV_60 $T=103960 204000 1 0 $X=103770 $Y=201040
X2895 VSS VDD 541 357 576 ICV_60 $T=103960 214880 1 0 $X=103770 $Y=211920
X2896 VSS VDD SCAN_IN<18> 749 767 ICV_60 $T=145820 78880 0 0 $X=145630 $Y=78640
X2897 VSS VDD 728 738 713 ICV_60 $T=145820 198560 0 0 $X=145630 $Y=198320
X2898 VSS VDD 821 818 762 ICV_60 $T=160080 19040 1 0 $X=159890 $Y=16080
X2899 VSS VDD 879 887 513 ICV_60 $T=173880 46240 0 0 $X=173690 $Y=46000
X2900 VSS VDD 881 888 802 ICV_60 $T=173880 84320 0 0 $X=173690 $Y=84080
X2901 VSS VDD 861 848 881 ICV_60 $T=173880 95200 0 0 $X=173690 $Y=94960
X2902 VSS VDD 919 927 926 ICV_60 $T=188140 89760 1 0 $X=187950 $Y=86800
X2903 VSS VDD SCAN_IN<3> 947 961 ICV_60 $T=188140 198560 1 0 $X=187950 $Y=195600
X2904 VSS VDD SCAN_IN<3> 823 948 ICV_60 $T=188140 209440 1 0 $X=187950 $Y=206480
X2905 VSS VDD 999 930 958 ICV_60 $T=201940 40800 0 0 $X=201750 $Y=40560
X2906 VSS VDD 308 315 257 ICV_61 $T=57040 127840 1 0 $X=56850 $Y=124880
X2907 VSS VDD 500 481 343 ICV_61 $T=94760 198560 1 0 $X=94570 $Y=195600
X2908 VSS VDD 714 735 725 ICV_61 $T=138460 35360 1 0 $X=138270 $Y=32400
X2909 VSS VDD 830 865 842 ICV_61 $T=176180 29920 1 0 $X=175990 $Y=26960
X2910 VSS VDD 900 913 876 ICV_61 $T=177100 127840 1 0 $X=176910 $Y=124880
X2911 VSS VDD 929 819 712 ICV_61 $T=189520 155040 1 0 $X=189330 $Y=152080
X2912 VSS VDD SCAN_IN<0> 929 991 ICV_61 $T=197800 160480 1 0 $X=197610 $Y=157520
X2913 VSS VDD 990 968 1010 ICV_61 $T=201480 225760 1 0 $X=201290 $Y=222800
X2914 VSS VDD 62 37 26 64 VDD 44 VSS sky130_fd_sc_hd__or4_4 $T=11960 89760 1 0 $X=11770 $Y=86800
X2915 VSS VDD 112 37 120 64 VDD 81 VSS sky130_fd_sc_hd__or4_4 $T=21160 89760 1 0 $X=20970 $Y=86800
X2916 VSS VDD 239 235 205 241 VDD 262 VSS sky130_fd_sc_hd__or4_4 $T=41860 73440 0 0 $X=41670 $Y=73200
X2917 VSS VDD 264 273 262 224 VDD 303 VSS sky130_fd_sc_hd__or4_4 $T=49220 51680 1 0 $X=49030 $Y=48720
X2918 VSS VDD 220 344 342 332 VDD 362 VSS sky130_fd_sc_hd__or4_4 $T=61640 68000 1 0 $X=61450 $Y=65040
X2919 VSS VDD 360 341 369 354 VDD 375 VSS sky130_fd_sc_hd__or4_4 $T=65320 73440 0 0 $X=65130 $Y=73200
X2920 VSS VDD 377 388 324 355 VDD 404 VSS sky130_fd_sc_hd__or4_4 $T=70380 133280 0 0 $X=70190 $Y=133040
X2921 VSS VDD 498 478 488 431 VDD 221 VSS sky130_fd_sc_hd__or4_4 $T=94300 127840 1 0 $X=94110 $Y=124880
X2922 VSS VDD 558 678 673 618 VDD 409 VSS sky130_fd_sc_hd__or4_4 $T=132020 155040 0 0 $X=131830 $Y=154800
X2923 VSS VDD 720 729 732 722 VDD 597 VSS sky130_fd_sc_hd__or4_4 $T=137080 111520 0 0 $X=136890 $Y=111280
X2924 VSS VDD 911 765 904 666 VDD 860 VSS sky130_fd_sc_hd__or4_4 $T=178480 62560 1 0 $X=178290 $Y=59600
X2925 VSS VDD 940 1003 977 987 VDD 898 VSS sky130_fd_sc_hd__or4_4 $T=201020 111520 1 0 $X=200830 $Y=108560
X2926 VSS 94 ICV_62 $T=17940 138720 1 0 $X=17750 $Y=135760
X2927 VSS 102 ICV_62 $T=17940 176800 1 0 $X=17750 $Y=173840
X2928 VSS 106 ICV_62 $T=17940 198560 1 0 $X=17750 $Y=195600
X2929 VSS 87 ICV_62 $T=17940 204000 1 0 $X=17750 $Y=201040
X2930 VSS 191 ICV_62 $T=31740 19040 0 0 $X=31550 $Y=18800
X2931 VSS 128 ICV_62 $T=31740 35360 0 0 $X=31550 $Y=35120
X2932 VSS 153 ICV_62 $T=31740 57120 0 0 $X=31550 $Y=56880
X2933 VSS 192 ICV_62 $T=31740 62560 0 0 $X=31550 $Y=62320
X2934 VSS 193 ICV_62 $T=31740 68000 0 0 $X=31550 $Y=67760
X2935 VSS 175 ICV_62 $T=31740 122400 0 0 $X=31550 $Y=122160
X2936 VSS 195 ICV_62 $T=31740 133280 0 0 $X=31550 $Y=133040
X2937 VSS 57 ICV_62 $T=31740 155040 0 0 $X=31550 $Y=154800
X2938 VSS 102 ICV_62 $T=31740 176800 0 0 $X=31550 $Y=176560
X2939 VSS 264 ICV_62 $T=46000 46240 1 0 $X=45810 $Y=43280
X2940 VSS 247 ICV_62 $T=46000 127840 1 0 $X=45810 $Y=124880
X2941 VSS 268 ICV_62 $T=46000 165920 1 0 $X=45810 $Y=162960
X2942 VSS 191 ICV_62 $T=59800 19040 0 0 $X=59610 $Y=18800
X2943 VSS 285 ICV_62 $T=59800 73440 0 0 $X=59610 $Y=73200
X2944 VSS 334 ICV_62 $T=59800 100640 0 0 $X=59610 $Y=100400
X2945 VSS 212 ICV_62 $T=59800 111520 0 0 $X=59610 $Y=111280
X2946 VSS 308 ICV_62 $T=59800 127840 0 0 $X=59610 $Y=127600
X2947 VSS 336 ICV_62 $T=59800 155040 0 0 $X=59610 $Y=154800
X2948 VSS 301 ICV_62 $T=59800 209440 0 0 $X=59610 $Y=209200
X2949 VSS 405 ICV_62 $T=74060 78880 1 0 $X=73870 $Y=75920
X2950 VSS CLK_IN ICV_62 $T=87860 13600 0 0 $X=87670 $Y=13360
X2951 VSS 326 ICV_62 $T=87860 100640 0 0 $X=87670 $Y=100400
X2952 VSS 190 ICV_62 $T=87860 182240 0 0 $X=87670 $Y=182000
X2953 VSS 464 ICV_62 $T=87860 214880 0 0 $X=87670 $Y=214640
X2954 VSS 464 ICV_62 $T=89240 225760 0 0 $X=89050 $Y=225520
X2955 VSS 538 ICV_62 $T=102120 176800 1 0 $X=101930 $Y=173840
X2956 VSS 506 ICV_62 $T=102120 182240 1 0 $X=101930 $Y=179280
X2957 VSS 541 ICV_62 $T=102120 209440 1 0 $X=101930 $Y=206480
X2958 VSS 614 ICV_62 $T=115920 78880 0 0 $X=115730 $Y=78640
X2959 VSS SCAN_IN<14> ICV_62 $T=115920 133280 0 0 $X=115730 $Y=133040
X2960 VSS SCAN_IN<16> ICV_62 $T=115920 138720 0 0 $X=115730 $Y=138480
X2961 VSS 549 ICV_62 $T=115920 160480 0 0 $X=115730 $Y=160240
X2962 VSS 618 ICV_62 $T=115920 165920 0 0 $X=115730 $Y=165680
X2963 VSS 620 ICV_62 $T=115920 193120 0 0 $X=115730 $Y=192880
X2964 VSS 321 ICV_62 $T=115920 204000 0 0 $X=115730 $Y=203760
X2965 VSS 290 ICV_62 $T=115920 220320 0 0 $X=115730 $Y=220080
X2966 VSS 393 ICV_62 $T=130180 84320 1 0 $X=129990 $Y=81360
X2967 VSS 661 ICV_62 $T=130180 127840 1 0 $X=129990 $Y=124880
X2968 VSS 697 ICV_62 $T=132020 13600 1 0 $X=131830 $Y=10640
X2969 VSS 755 ICV_62 $T=143980 51680 0 0 $X=143790 $Y=51440
X2970 VSS 758 ICV_62 $T=143980 127840 0 0 $X=143790 $Y=127600
X2971 VSS 761 ICV_62 $T=143980 165920 0 0 $X=143790 $Y=165680
X2972 VSS 803 ICV_62 $T=158240 68000 1 0 $X=158050 $Y=65040
X2973 VSS 703 ICV_62 $T=158240 84320 1 0 $X=158050 $Y=81360
X2974 VSS 811 ICV_62 $T=158240 95200 1 0 $X=158050 $Y=92240
X2975 VSS 20 ICV_62 $T=158240 165920 1 0 $X=158050 $Y=162960
X2976 VSS 890 ICV_62 $T=172040 29920 0 0 $X=171850 $Y=29680
X2977 VSS 888 ICV_62 $T=172040 78880 0 0 $X=171850 $Y=78640
X2978 VSS 892 ICV_62 $T=172040 116960 0 0 $X=171850 $Y=116720
X2979 VSS 846 ICV_62 $T=172040 138720 0 0 $X=171850 $Y=138480
X2980 VSS 896 ICV_62 $T=172040 182240 0 0 $X=171850 $Y=182000
X2981 VSS 507 ICV_62 $T=172040 204000 0 0 $X=171850 $Y=203760
X2982 VSS 855 ICV_62 $T=172040 220320 0 0 $X=171850 $Y=220080
X2983 VSS 944 ICV_62 $T=186300 100640 1 0 $X=186110 $Y=97680
X2984 VSS 946 ICV_62 $T=186300 182240 1 0 $X=186110 $Y=179280
X2985 VSS 999 ICV_62 $T=200100 35360 0 0 $X=199910 $Y=35120
X2986 VSS 784 ICV_62 $T=200100 57120 0 0 $X=199910 $Y=56880
X2987 VSS 1001 ICV_62 $T=200100 73440 0 0 $X=199910 $Y=73200
X2988 VSS 977 ICV_62 $T=200100 106080 0 0 $X=199910 $Y=105840
X2989 VSS 1003 ICV_62 $T=200100 122400 0 0 $X=199910 $Y=122160
X2990 VSS 158 ICV_62 $T=200100 127840 0 0 $X=199910 $Y=127600
X2991 VSS 984 ICV_62 $T=200100 171360 0 0 $X=199910 $Y=171120
X2992 VSS 957 ICV_62 $T=200100 214880 0 0 $X=199910 $Y=214640
X2993 VSS VDD 106 ICV_63 $T=17940 193120 1 0 $X=17750 $Y=190160
X2994 VSS VDD 187 ICV_63 $T=31740 138720 0 0 $X=31550 $Y=138480
X2995 VSS VDD 406 ICV_63 $T=74060 133280 1 0 $X=73870 $Y=130320
X2996 VSS VDD 407 ICV_63 $T=74060 155040 1 0 $X=73870 $Y=152080
X2997 VSS VDD 441 ICV_63 $T=87860 160480 0 0 $X=87670 $Y=160240
X2998 VSS VDD 540 ICV_63 $T=102120 193120 1 0 $X=101930 $Y=190160
X2999 VSS VDD 591 ICV_63 $T=115920 35360 0 0 $X=115730 $Y=35120
X3000 VSS VDD 644 ICV_63 $T=143980 106080 0 0 $X=143790 $Y=105840
X3001 VSS VDD 796 ICV_63 $T=158240 57120 1 0 $X=158050 $Y=54160
X3002 VSS VDD 961 ICV_63 $T=200100 187680 0 0 $X=199910 $Y=187440
X3003 VSS VDD 24 73 25 VDD 42 VSS sky130_fd_sc_hd__a21o_4 $T=7820 62560 0 0 $X=7630 $Y=62320
X3004 VSS VDD 69 SCAN_IN<9> 33 VDD 39 VSS sky130_fd_sc_hd__a21o_4 $T=8740 165920 0 0 $X=8550 $Y=165680
X3005 VSS VDD 150 166 125 VDD 78 VSS sky130_fd_sc_hd__a21o_4 $T=22540 193120 1 0 $X=22350 $Y=190160
X3006 VSS VDD 79 138 127 VDD 151 VSS sky130_fd_sc_hd__a21o_4 $T=23460 214880 0 0 $X=23270 $Y=214640
X3007 VSS VDD 150 166 144 VDD 126 VSS sky130_fd_sc_hd__a21o_4 $T=23920 198560 1 0 $X=23730 $Y=195600
X3008 VSS VDD 217 214 194 VDD 159 VSS sky130_fd_sc_hd__a21o_4 $T=38640 111520 1 0 $X=38450 $Y=108560
X3009 VSS VDD 132 286 271 VDD 282 VSS sky130_fd_sc_hd__a21o_4 $T=49220 182240 1 0 $X=49030 $Y=179280
X3010 VSS VDD 150 166 340 VDD 314 VSS sky130_fd_sc_hd__a21o_4 $T=63020 198560 0 0 $X=62830 $Y=198320
X3011 VSS VDD 397 391 383 VDD 376 VSS sky130_fd_sc_hd__a21o_4 $T=74520 29920 0 0 $X=74330 $Y=29680
X3012 VSS VDD 425 SCAN_IN<7> 331 VDD 429 VSS sky130_fd_sc_hd__a21o_4 $T=78660 155040 1 0 $X=78470 $Y=152080
X3013 VSS VDD 338 433 441 VDD 415 VSS sky130_fd_sc_hd__a21o_4 $T=81420 182240 1 0 $X=81230 $Y=179280
X3014 VSS VDD 401 58 451 VDD 459 VSS sky130_fd_sc_hd__a21o_4 $T=85560 198560 1 0 $X=85370 $Y=195600
X3015 VSS VDD 502 513 519 VDD 453 VSS sky130_fd_sc_hd__a21o_4 $T=98900 46240 0 0 $X=98710 $Y=46000
X3016 VSS VDD 520 521 417 VDD 524 VSS sky130_fd_sc_hd__a21o_4 $T=98900 73440 0 0 $X=98710 $Y=73200
X3017 VSS VDD 528 512 506 VDD 479 VSS sky130_fd_sc_hd__a21o_4 $T=98900 165920 0 0 $X=98710 $Y=165680
X3018 VSS VDD 401 557 145 VDD 543 VSS sky130_fd_sc_hd__a21o_4 $T=101660 198560 0 0 $X=101470 $Y=198320
X3019 VSS VDD 520 521 452 VDD 564 VSS sky130_fd_sc_hd__a21o_4 $T=105340 51680 1 0 $X=105150 $Y=48720
X3020 VSS VDD 491 535 547 VDD 557 VSS sky130_fd_sc_hd__a21o_4 $T=105340 204000 0 0 $X=105150 $Y=203760
X3021 VSS VDD 499 550 590 VDD 484 VSS sky130_fd_sc_hd__a21o_4 $T=105800 176800 0 0 $X=105610 $Y=176560
X3022 VSS VDD 533 SCAN_IN<9> 525 VDD 586 VSS sky130_fd_sc_hd__a21o_4 $T=108100 24480 1 0 $X=107910 $Y=21520
X3023 VSS VDD 401 58 515 VDD 602 VSS sky130_fd_sc_hd__a21o_4 $T=111780 204000 1 0 $X=111590 $Y=201040
X3024 VSS VDD 643 607 534 VDD 638 VSS sky130_fd_sc_hd__a21o_4 $T=119140 57120 0 0 $X=118950 $Y=56880
X3025 VSS VDD 631 674 676 VDD 694 VSS sky130_fd_sc_hd__a21o_4 $T=130180 29920 0 0 $X=129990 $Y=29680
X3026 VSS VDD 646 728 738 VDD 579 VSS sky130_fd_sc_hd__a21o_4 $T=135240 204000 1 0 $X=135050 $Y=201040
X3027 VSS VDD 520 521 443 VDD 782 VSS sky130_fd_sc_hd__a21o_4 $T=150880 51680 0 0 $X=150690 $Y=51440
X3028 VSS VDD 787 596 503 VDD 825 VSS sky130_fd_sc_hd__a21o_4 $T=160540 84320 0 0 $X=160350 $Y=84080
X3029 VSS VDD 787 596 530 VDD 827 VSS sky130_fd_sc_hd__a21o_4 $T=160540 111520 0 0 $X=160350 $Y=111280
X3030 VSS VDD 787 826 608 VDD 811 VSS sky130_fd_sc_hd__a21o_4 $T=161460 95200 1 0 $X=161270 $Y=92240
X3031 VSS VDD 696 786 SCAN_IN<0> VDD 837 VSS sky130_fd_sc_hd__a21o_4 $T=162380 204000 0 0 $X=162190 $Y=203760
X3032 VSS VDD 867 861 848 VDD 826 VSS sky130_fd_sc_hd__a21o_4 $T=169740 95200 1 0 $X=169550 $Y=92240
X3033 VSS VDD 815 885 875 VDD 454 VSS sky130_fd_sc_hd__a21o_4 $T=171120 57120 1 0 $X=170930 $Y=54160
X3034 VSS VDD 853 SCAN_IN<7> 887 VDD 918 VSS sky130_fd_sc_hd__a21o_4 $T=178020 19040 1 0 $X=177830 $Y=16080
X3035 VSS VDD 921 919 927 VDD 511 VSS sky130_fd_sc_hd__a21o_4 $T=180780 89760 0 0 $X=180590 $Y=89520
X3036 VSS VDD 909 712 928 VDD 592 VSS sky130_fd_sc_hd__a21o_4 $T=181240 116960 0 0 $X=181050 $Y=116720
X3037 VSS VDD 901 SCAN_IN<1> 855 VDD 957 VSS sky130_fd_sc_hd__a21o_4 $T=189060 220320 0 0 $X=188870 $Y=220080
X3038 VSS VDD 944 774 848 VDD 922 VSS sky130_fd_sc_hd__a21o_4 $T=189520 106080 1 0 $X=189330 $Y=103120
X3039 VSS VDD 964 963 912 VDD 955 VSS sky130_fd_sc_hd__a21o_4 $T=190900 68000 1 0 $X=190710 $Y=65040
X3040 VSS VDD 978 991 998 VDD 1005 VSS sky130_fd_sc_hd__a21o_4 $T=199640 165920 1 0 $X=199450 $Y=162960
X3041 VSS VDD 25 63 ICV_64 $T=7820 68000 1 0 $X=7630 $Y=65040
X3042 VSS VDD 27 64 ICV_64 $T=7820 95200 0 0 $X=7630 $Y=94960
X3043 VSS VDD 68 105 ICV_64 $T=17020 155040 0 0 $X=16830 $Y=154800
X3044 VSS VDD 88 133 ICV_64 $T=21160 24480 0 0 $X=20970 $Y=24240
X3045 VSS VDD 172 172 ICV_64 $T=29440 89760 0 0 $X=29250 $Y=89520
X3046 VSS VDD 184 231 ICV_64 $T=37260 204000 0 0 $X=37070 $Y=203760
X3047 VSS VDD SCAN_IN<20> 188 ICV_64 $T=40480 138720 0 0 $X=40290 $Y=138480
X3048 VSS VDD 302 312 ICV_64 $T=52440 29920 1 0 $X=52250 $Y=26960
X3049 VSS VDD 147 390 ICV_64 $T=68080 19040 0 0 $X=67890 $Y=18800
X3050 VSS VDD 626 642 ICV_64 $T=118220 204000 1 0 $X=118030 $Y=201040
X3051 VSS VDD 770 795 ICV_64 $T=151340 198560 0 0 $X=151150 $Y=198320
X3052 VSS VDD 755 808 ICV_64 $T=160540 133280 0 0 $X=160350 $Y=133040
X3053 VSS VDD 418 887 ICV_64 $T=169740 13600 0 0 $X=169550 $Y=13360
X3054 VSS VDD 769 769 ICV_64 $T=169740 149600 0 0 $X=169550 $Y=149360
X3055 VSS VDD 618 895 ICV_64 $T=169740 176800 0 0 $X=169550 $Y=176560
X3056 VSS VDD 881 574 ICV_64 $T=172040 84320 1 0 $X=171850 $Y=81360
X3057 VSS VDD 842 935 ICV_64 $T=192280 29920 0 0 $X=192090 $Y=29680
X3058 VSS VDD 940 985 ICV_64 $T=198720 133280 1 0 $X=198530 $Y=130320
X3059 VSS 26 44 ICV_65 $T=16100 95200 1 0 $X=15910 $Y=92240
X3060 VSS 39 103 ICV_65 $T=16100 165920 1 0 $X=15910 $Y=162960
X3061 VSS 205 267 ICV_65 $T=44160 78880 1 0 $X=43970 $Y=75920
X3062 VSS 326 334 ICV_65 $T=57960 95200 0 0 $X=57770 $Y=94960
X3063 VSS 321 248 ICV_65 $T=57960 171360 0 0 $X=57770 $Y=171120
X3064 VSS 189 339 ICV_65 $T=57960 193120 0 0 $X=57770 $Y=192880
X3065 VSS 452 448 ICV_65 $T=86020 57120 0 0 $X=85830 $Y=56880
X3066 VSS 456 20 ICV_65 $T=86020 155040 0 0 $X=85830 $Y=154800
X3067 VSS 321 469 ICV_65 $T=86020 187680 0 0 $X=85830 $Y=187440
X3068 VSS 295 537 ICV_65 $T=100280 149600 1 0 $X=100090 $Y=146640
X3069 VSS 145 539 ICV_65 $T=100280 187680 1 0 $X=100090 $Y=184720
X3070 VSS 554 533 ICV_65 $T=114080 19040 0 0 $X=113890 $Y=18800
X3071 VSS 608 525 ICV_65 $T=114080 29920 0 0 $X=113890 $Y=29680
X3072 VSS 534 534 ICV_65 $T=114080 57120 0 0 $X=113890 $Y=56880
X3073 VSS 575 615 ICV_65 $T=114080 116960 0 0 $X=113890 $Y=116720
X3074 VSS 458 617 ICV_65 $T=114080 144160 0 0 $X=113890 $Y=143920
X3075 VSS 456 689 ICV_65 $T=128340 78880 1 0 $X=128150 $Y=75920
X3076 VSS 748 628 ICV_65 $T=142140 35360 0 0 $X=141950 $Y=35120
X3077 VSS 749 SCAN_IN<18> ICV_65 $T=142140 84320 0 0 $X=141950 $Y=84080
X3078 VSS 422 756 ICV_65 $T=142140 95200 0 0 $X=141950 $Y=94960
X3079 VSS SCAN_IN<13> 759 ICV_65 $T=142140 144160 0 0 $X=141950 $Y=143920
X3080 VSS 751 590 ICV_65 $T=142140 176800 0 0 $X=141950 $Y=176560
X3081 VSS 738 680 ICV_65 $T=142140 182240 0 0 $X=141950 $Y=182000
X3082 VSS 738 680 ICV_65 $T=142140 187680 0 0 $X=141950 $Y=187440
X3083 VSS 634 747 ICV_65 $T=142140 220320 0 0 $X=141950 $Y=220080
X3084 VSS 878 878 ICV_65 $T=170200 19040 0 0 $X=170010 $Y=18800
X3085 VSS 938 948 ICV_65 $T=184460 214880 1 0 $X=184270 $Y=211920
X3086 VSS 995 996 ICV_65 $T=198260 84320 0 0 $X=198070 $Y=84080
X3087 VSS 996 976 ICV_65 $T=198260 95200 0 0 $X=198070 $Y=94960
X3088 VSS VDD 86 ICV_66 $T=16100 89760 1 0 $X=15910 $Y=86800
X3089 VSS VDD 408 ICV_66 $T=72220 171360 1 0 $X=72030 $Y=168400
X3090 VSS VDD 524 ICV_66 $T=100280 68000 1 0 $X=100090 $Y=65040
X3091 VSS VDD 607 ICV_66 $T=114080 62560 0 0 $X=113890 $Y=62320
X3092 VSS VDD 631 ICV_66 $T=128340 35360 1 0 $X=128150 $Y=32400
X3093 VSS VDD 757 ICV_66 $T=142140 122400 0 0 $X=141950 $Y=122160
X3094 VSS VDD 703 ICV_66 $T=156400 100640 1 0 $X=156210 $Y=97680
X3095 VSS VDD 865 ICV_66 $T=170200 35360 0 0 $X=170010 $Y=35120
X3096 VSS VDD 20 ICV_66 $T=198260 46240 0 0 $X=198070 $Y=46000
X3097 VSS VDD 124 259 238 ICV_67 $T=42320 19040 0 0 $X=42130 $Y=18800
X3098 VSS VDD 171 277 276 ICV_67 $T=45080 78880 0 0 $X=44890 $Y=78640
X3099 VSS VDD 273 318 307 ICV_67 $T=54740 46240 0 0 $X=54550 $Y=46000
X3100 VSS VDD 351 128 373 ICV_67 $T=63020 46240 0 0 $X=62830 $Y=46000
X3101 VSS VDD 655 253 666 ICV_67 $T=126960 19040 0 0 $X=126770 $Y=18800
X3102 VSS VDD SCAN_IN<13> 721 757 ICV_67 $T=147200 133280 0 0 $X=147010 $Y=133040
X3103 VSS VDD 744 802 810 ICV_67 $T=153640 57120 0 0 $X=153450 $Y=56880
X3104 VSS VDD 957 968 990 ICV_67 $T=195500 220320 0 0 $X=195310 $Y=220080
X3105 VSS VDD 105 132 87 59 143 VDD 125 VSS sky130_fd_sc_hd__a32o_4 $T=22080 182240 0 0 $X=21890 $Y=182000
X3106 VSS VDD 195 221 228 SCAN_IN<21> 95 VDD 176 VSS sky130_fd_sc_hd__a32o_4 $T=36340 138720 1 0 $X=36150 $Y=135760
X3107 VSS VDD 186 236 243 246 192 VDD 223 VSS sky130_fd_sc_hd__a32o_4 $T=38180 62560 0 0 $X=37990 $Y=62320
X3108 VSS VDD 260 250 232 191 238 VDD 62 VSS sky130_fd_sc_hd__a32o_4 $T=43240 29920 0 0 $X=43050 $Y=29680
X3109 VSS VDD 244 269 268 231 256 VDD 131 VSS sky130_fd_sc_hd__a32o_4 $T=46000 165920 0 0 $X=45810 $Y=165680
X3110 VSS VDD 510 502 489 529 501 VDD 417 VSS sky130_fd_sc_hd__a32o_4 $T=97980 51680 0 0 $X=97790 $Y=51440
X3111 VSS VDD 582 581 401 553 544 VDD 563 VSS sky130_fd_sc_hd__a32o_4 $T=106260 220320 1 0 $X=106070 $Y=217360
X3112 VSS VDD 599 597 588 SCAN_IN<21> 573 VDD 566 VSS sky130_fd_sc_hd__a32o_4 $T=111320 106080 1 0 $X=111130 $Y=103120
X3113 VSS VDD 777 793 787 794 800 VDD 792 VSS sky130_fd_sc_hd__a32o_4 $T=152720 155040 0 0 $X=152530 $Y=154800
X3114 VSS VDD 842 756 810 788 830 VDD 773 VSS sky130_fd_sc_hd__a32o_4 $T=161920 35360 1 0 $X=161730 $Y=32400
X3115 VSS VDD 948 SCAN_IN<2> 795 823 SCAN_IN<3> VDD 938 VSS sky130_fd_sc_hd__a32o_4 $T=187220 209440 0 0 $X=187030 $Y=209200
X3116 VSS VDD 916 SCAN_IN<4> 801 532 SCAN_IN<5> VDD 931 VSS sky130_fd_sc_hd__a32o_4 $T=189520 171360 1 0 $X=189330 $Y=168400
X3117 VSS VDD 950 SCAN_IN<4> 927 956 SCAN_IN<5> VDD 970 VSS sky130_fd_sc_hd__a32o_4 $T=194120 84320 1 0 $X=193930 $Y=81360
X3118 VSS VDD 961 SCAN_IN<2> 960 913 SCAN_IN<3> VDD 979 VSS sky130_fd_sc_hd__a32o_4 $T=195500 198560 1 0 $X=195310 $Y=195600
X3119 VSS VDD 22 19 77 ICV_68 $T=7820 40800 0 0 $X=7630 $Y=40560
X3120 VSS VDD 161 206 206 ICV_68 $T=36340 198560 0 0 $X=36150 $Y=198320
X3121 VSS VDD 298 288 317 ICV_68 $T=51520 24480 1 0 $X=51330 $Y=21520
X3122 VSS VDD 422 439 20 ICV_68 $T=83260 116960 0 0 $X=83070 $Y=116720
X3123 VSS VDD 604 522 522 ICV_68 $T=119140 46240 0 0 $X=118950 $Y=46000
X3124 VSS VDD 734 437 495 ICV_68 $T=139380 214880 0 0 $X=139190 $Y=214640
X3125 VSS VDD 521 859 893 ICV_68 $T=167440 122400 0 0 $X=167250 $Y=122160
X3126 VSS VDD 532 916 984 ICV_68 $T=195500 165920 0 0 $X=195310 $Y=165680
X3127 VSS VDD 232 ICV_69 $T=38180 35360 0 0 $X=37990 $Y=35120
X3128 VSS VDD 333 ICV_69 $T=56120 57120 1 0 $X=55930 $Y=54160
X3129 VSS VDD 326 ICV_69 $T=79120 106080 0 0 $X=78930 $Y=105840
X3130 VSS VDD 463 ICV_69 $T=83260 220320 1 0 $X=83070 $Y=217360
X3131 VSS VDD 666 ICV_69 $T=151800 19040 0 0 $X=151610 $Y=18800
X3132 VSS VDD 896 ICV_69 $T=171580 187680 1 0 $X=171390 $Y=184720
X3133 VSS VDD 650 ICV_69 $T=191360 68000 0 0 $X=191170 $Y=67760
X3134 VSS VDD 997 ICV_69 $T=195040 127840 1 0 $X=194850 $Y=124880
X3135 VSS VDD 159 ICV_70 $T=25760 100640 1 0 $X=25570 $Y=97680
X3136 VSS VDD 224 ICV_70 $T=37720 51680 0 0 $X=37530 $Y=51440
X3137 VSS VDD 289 ICV_70 $T=48300 68000 1 0 $X=48110 $Y=65040
X3138 VSS VDD 272 ICV_70 $T=51060 204000 0 0 $X=50870 $Y=203760
X3139 VSS VDD 189 ICV_70 $T=116840 193120 1 0 $X=116650 $Y=190160
X3140 VSS VDD 237 ICV_70 $T=122820 193120 1 0 $X=122630 $Y=190160
X3141 VSS VDD 879 ICV_70 $T=172960 46240 1 0 $X=172770 $Y=43280
X3142 VSS VDD 977 ICV_70 $T=194120 106080 0 0 $X=193930 $Y=105840
X3143 VSS VDD 85 85 168 117 ICV_71 $T=24840 40800 0 0 $X=24650 $Y=40560
X3144 VSS VDD 229 229 179 234 ICV_71 $T=39100 84320 0 0 $X=38910 $Y=84080
X3145 VSS VDD 257 257 247 175 ICV_71 $T=46460 127840 0 0 $X=46270 $Y=127600
X3146 VSS VDD 283 297 310 283 ICV_71 $T=51520 225760 1 0 $X=51330 $Y=222800
X3147 VSS VDD 43 43 275 323 ICV_71 $T=52900 68000 0 0 $X=52710 $Y=67760
X3148 VSS VDD 297 343 349 297 ICV_71 $T=60260 220320 1 0 $X=60070 $Y=217360
X3149 VSS VDD 357 398 357 399 ICV_71 $T=70380 209440 0 0 $X=70190 $Y=209200
X3150 VSS VDD 441 433 441 353 ICV_71 $T=80960 176800 0 0 $X=80770 $Y=176560
X3151 VSS VDD 493 493 525 501 ICV_71 $T=97980 35360 0 0 $X=97790 $Y=35120
X3152 VSS VDD 549 561 568 526 ICV_71 $T=103960 149600 0 0 $X=103770 $Y=149360
X3153 VSS VDD 590 550 590 538 ICV_71 $T=109480 182240 1 0 $X=109290 $Y=179280
X3154 VSS VDD 692 692 641 535 ICV_71 $T=130180 209440 0 0 $X=129990 $Y=209200
X3155 VSS VDD 784 SCAN_IN<16> 784 710 ICV_71 $T=150420 100640 0 0 $X=150230 $Y=100400
X3156 VSS VDD 790 859 521 816 ICV_71 $T=165600 127840 1 0 $X=165410 $Y=124880
X3157 VSS VDD 20 926 912 885 ICV_71 $T=179400 78880 1 0 $X=179210 $Y=75920
X3158 VSS VDD 928 712 928 923 ICV_71 $T=184460 122400 0 0 $X=184270 $Y=122160
X3159 VSS VDD SCAN_IN<4> SCAN_IN<5> 956 950 ICV_71 $T=193200 78880 0 0 $X=193010 $Y=78640
X3160 VSS VDD 133 147 116 147 ICV_72 $T=22540 19040 0 0 $X=22350 $Y=18800
X3161 VSS VDD 312 84 302 84 ICV_72 $T=51060 29920 0 0 $X=50870 $Y=29680
X3162 VSS VDD 513 519 493 519 ICV_72 $T=99360 40800 0 0 $X=99170 $Y=40560
X3163 VSS VDD 663 166 654 654 ICV_72 $T=120520 225760 1 0 $X=120330 $Y=222800
X3164 VSS VDD 902 519 884 519 ICV_72 $T=181240 35360 0 0 $X=181050 $Y=35120
X3165 VSS VDD 923 913 919 913 ICV_72 $T=186760 116960 0 0 $X=186570 $Y=116720
X3166 VSS VDD SCAN_IN<5> 532 916 532 ICV_72 $T=188140 171360 0 0 $X=187950 $Y=171120
X3167 VSS VDD 958 902 670 958 ICV_72 $T=190440 51680 0 0 $X=190250 $Y=51440
X3168 VSS VDD 723 721 989 721 ICV_72 $T=191360 133280 0 0 $X=191170 $Y=133040
X3169 VSS VDD 32 57 33 ICV_73 $T=7820 171360 1 0 $X=7630 $Y=168400
X3170 VSS VDD 152 64 140 ICV_73 $T=23460 100640 0 0 $X=23270 $Y=100400
X3171 VSS VDD 173 59 176 ICV_73 $T=28060 176800 1 0 $X=27870 $Y=173840
X3172 VSS VDD 234 243 235 ICV_73 $T=40020 78880 1 0 $X=39830 $Y=75920
X3173 VSS VDD 258 127 231 ICV_73 $T=45080 193120 0 0 $X=44890 $Y=192880
X3174 VSS VDD 326 509 17 ICV_73 $T=93380 100640 0 0 $X=93190 $Y=100400
X3175 VSS VDD 656 664 664 ICV_73 $T=124200 95200 0 0 $X=124010 $Y=94960
X3176 VSS VDD 744 790 622 ICV_73 $T=149500 57120 0 0 $X=149310 $Y=56880
X3177 VSS VDD 801 590 779 ICV_73 $T=154560 176800 0 0 $X=154370 $Y=176560
X3178 VSS VDD 745 608 745 ICV_73 $T=155480 84320 0 0 $X=155290 $Y=84080
X3179 VSS VDD 945 927 945 ICV_73 $T=190900 106080 0 0 $X=190710 $Y=105840
X3180 VSS VDD 109 137 158 102 113 100 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=21160 138720 1 0 $X=20970 $Y=135760
X3181 VSS VDD 109 93 158 136 175 156 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=24380 133280 1 0 $X=24190 $Y=130320
X3182 VSS VDD 109 549 466 537 471 569 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=105340 155040 1 0 $X=105150 $Y=152080
X3183 VSS VDD 548 346 536 565 562 567 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=105800 95200 1 0 $X=105610 $Y=92240
X3184 VSS VDD 937 962 954 875 930 748 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=189520 40800 1 0 $X=189330 $Y=37840
X3185 VSS VDD BB_IN 13 ICV_74 $T=7820 138720 0 0 $X=7630 $Y=138480
X3186 VSS VDD 59 58 ICV_74 $T=9660 198560 0 0 $X=9470 $Y=198320
X3187 VSS VDD 62 27 ICV_74 $T=12880 100640 1 0 $X=12690 $Y=97680
X3188 VSS VDD 43 55 ICV_74 $T=21160 73440 0 0 $X=20970 $Y=73200
X3189 VSS VDD 121 160 ICV_74 $T=24840 122400 0 0 $X=24650 $Y=122160
X3190 VSS VDD 118 131 ICV_74 $T=26220 165920 0 0 $X=26030 $Y=165680
X3191 VSS VDD 225 245 ICV_74 $T=40480 204000 1 0 $X=40290 $Y=201040
X3192 VSS VDD 267 242 ICV_74 $T=49220 89760 1 0 $X=49030 $Y=86800
X3193 VSS VDD 379 392 ICV_74 $T=69000 62560 1 0 $X=68810 $Y=59600
X3194 VSS VDD 290 483 ICV_74 $T=95220 214880 0 0 $X=95030 $Y=214640
X3195 VSS VDD 481 500 ICV_74 $T=97060 193120 0 0 $X=96870 $Y=192880
X3196 VSS VDD 598 629 ICV_74 $T=119140 78880 0 0 $X=118950 $Y=78640
X3197 VSS VDD 598 562 ICV_74 $T=123280 84320 1 0 $X=123090 $Y=81360
X3198 VSS VDD 576 166 ICV_74 $T=125120 220320 1 0 $X=124930 $Y=217360
X3199 VSS VDD 787 608 ICV_74 $T=161460 89760 0 0 $X=161270 $Y=89520
X3200 VSS VDD 830 771 ICV_74 $T=162840 40800 1 0 $X=162650 $Y=37840
X3201 VSS VDD 804 836 ICV_74 $T=163760 176800 1 0 $X=163570 $Y=173840
X3202 VSS VDD 903 903 ICV_74 $T=175260 176800 1 0 $X=175070 $Y=173840
X3203 VSS VDD 928 909 ICV_74 $T=181240 122400 1 0 $X=181050 $Y=119440
X3204 VSS VDD 929 819 ICV_74 $T=188600 149600 0 0 $X=188410 $Y=149360
X3205 VSS VDD 211 172 179 229 199 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=35420 89760 1 0 $X=35230 $Y=86800
X3206 VSS VDD 410 378 339 364 408 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=77280 171360 1 0 $X=77090 $Y=168400
X3207 VSS VDD 340 448 458 443 435 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=84640 57120 1 0 $X=84450 $Y=54160
X3208 VSS VDD 479 482 441 476 319 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=89700 165920 1 0 $X=89510 $Y=162960
X3209 VSS VDD 144 448 458 452 445 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=91080 57120 0 0 $X=90890 $Y=56880
X3210 VSS VDD 451 448 458 503 450 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=92920 84320 0 0 $X=92730 $Y=84080
X3211 VSS VDD 515 448 393 530 497 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=99360 111520 0 0 $X=99170 $Y=111280
X3212 VSS VDD 836 568 337 804 840 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=161920 182240 1 0 $X=161730 $Y=179280
X3213 VSS VDD 922 934 888 771 937 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=183540 95200 0 0 $X=183350 $Y=94960
X3214 VSS VDD 955 959 875 784 906 VDD VSS sky130_fd_sc_hd__a22oi_4 $T=188600 57120 0 0 $X=188410 $Y=56880
X3215 VSS VDD ICV_75 $T=19780 62560 1 0 $X=19590 $Y=59600
X3216 VSS VDD ICV_75 $T=19780 68000 1 0 $X=19590 $Y=65040
X3217 VSS VDD ICV_75 $T=19780 100640 1 0 $X=19590 $Y=97680
X3218 VSS VDD ICV_75 $T=19780 155040 1 0 $X=19590 $Y=152080
X3219 VSS VDD ICV_75 $T=33580 95200 0 0 $X=33390 $Y=94960
X3220 VSS VDD ICV_75 $T=61640 89760 0 0 $X=61450 $Y=89520
X3221 VSS VDD ICV_75 $T=61640 116960 0 0 $X=61450 $Y=116720
X3222 VSS VDD ICV_75 $T=89700 29920 0 0 $X=89510 $Y=29680
X3223 VSS VDD ICV_75 $T=117760 13600 0 0 $X=117570 $Y=13360
X3224 VSS VDD ICV_75 $T=117760 24480 0 0 $X=117570 $Y=24240
X3225 VSS VDD ICV_75 $T=117760 95200 0 0 $X=117570 $Y=94960
X3226 VSS VDD ICV_75 $T=132020 122400 1 0 $X=131830 $Y=119440
X3227 VSS VDD ICV_75 $T=132020 171360 1 0 $X=131830 $Y=168400
X3228 VSS VDD ICV_75 $T=132020 176800 1 0 $X=131830 $Y=173840
X3229 VSS VDD ICV_75 $T=145820 19040 0 0 $X=145630 $Y=18800
X3230 VSS VDD ICV_75 $T=145820 24480 0 0 $X=145630 $Y=24240
X3231 VSS VDD ICV_75 $T=145820 111520 0 0 $X=145630 $Y=111280
X3232 VSS VDD ICV_75 $T=160080 122400 1 0 $X=159890 $Y=119440
X3233 VSS VDD ICV_75 $T=160080 160480 1 0 $X=159890 $Y=157520
X3234 VSS VDD ICV_75 $T=160080 171360 1 0 $X=159890 $Y=168400
X3235 VSS VDD ICV_75 $T=160080 225760 1 0 $X=159890 $Y=222800
X3236 VSS VDD ICV_75 $T=188140 19040 1 0 $X=187950 $Y=16080
X3237 VSS VDD ICV_75 $T=188140 111520 1 0 $X=187950 $Y=108560
X3238 VSS 147 139 170 ICV_76 $T=28060 13600 0 0 $X=27870 $Y=13360
X3239 VSS 157 168 20 ICV_76 $T=28060 46240 0 0 $X=27870 $Y=46000
X3240 VSS 318 307 307 ICV_76 $T=56120 51680 0 0 $X=55930 $Y=51440
X3241 VSS 282 453 466 ICV_76 $T=84180 73440 0 0 $X=83990 $Y=73200
X3242 VSS 20 450 466 ICV_76 $T=84180 78880 0 0 $X=83990 $Y=78640
X3243 VSS 506 512 528 ICV_76 $T=98440 165920 1 0 $X=98250 $Y=162960
X3244 VSS 740 551 676 ICV_76 $T=140300 40800 0 0 $X=140110 $Y=40560
X3245 VSS 741 325 760 ICV_76 $T=140300 160480 0 0 $X=140110 $Y=160240
X3246 VSS 783 614 730 ICV_76 $T=154560 78880 1 0 $X=154370 $Y=75920
X3247 VSS 863 SCAN_IN<0> 747 ICV_76 $T=168360 214880 0 0 $X=168170 $Y=214640
X3248 VSS 864 918 918 ICV_76 $T=185380 13600 1 0 $X=185190 $Y=10640
X3249 VSS VDD 16 51 20 VDD 105 VSS sky130_fd_sc_hd__dfstp_4 $T=7820 182240 0 0 $X=7630 $Y=182000
X3250 VSS VDD 16 52 20 VDD 33 VSS sky130_fd_sc_hd__dfstp_4 $T=7820 204000 0 0 $X=7630 $Y=203760
X3251 VSS VDD 16 183 20 VDD 249 VSS sky130_fd_sc_hd__dfstp_4 $T=32660 225760 1 0 $X=32470 $Y=222800
X3252 VSS VDD 212 233 20 VDD 194 VSS sky130_fd_sc_hd__dfstp_4 $T=39560 116960 0 0 $X=39370 $Y=116720
X3253 VSS VDD 212 296 20 VDD 214 VSS sky130_fd_sc_hd__dfstp_4 $T=49680 111520 1 0 $X=49490 $Y=108560
X3254 VSS VDD 16 311 20 VDD 331 VSS sky130_fd_sc_hd__dfstp_4 $T=52440 193120 1 0 $X=52250 $Y=190160
X3255 VSS VDD 416 427 20 VDD 275 VSS sky130_fd_sc_hd__dfstp_4 $T=77280 73440 1 0 $X=77090 $Y=70480
X3256 VSS VDD 16 411 20 VDD 441 VSS sky130_fd_sc_hd__dfstp_4 $T=77280 204000 1 0 $X=77090 $Y=201040
X3257 VSS VDD 416 434 20 VDD 412 VSS sky130_fd_sc_hd__dfstp_4 $T=78200 40800 1 0 $X=78010 $Y=37840
X3258 VSS VDD 416 435 20 VDD 330 VSS sky130_fd_sc_hd__dfstp_4 $T=78660 62560 1 0 $X=78470 $Y=59600
X3259 VSS VDD 416 440 20 VDD 373 VSS sky130_fd_sc_hd__dfstp_4 $T=79580 68000 1 0 $X=79390 $Y=65040
X3260 VSS VDD 416 445 20 VDD 383 VSS sky130_fd_sc_hd__dfstp_4 $T=81880 46240 1 0 $X=81690 $Y=43280
X3261 VSS VDD 416 450 20 VDD 276 VSS sky130_fd_sc_hd__dfstp_4 $T=84180 84320 1 0 $X=83990 $Y=81360
X3262 VSS VDD 416 455 20 VDD 266 VSS sky130_fd_sc_hd__dfstp_4 $T=84640 95200 1 0 $X=84450 $Y=92240
X3263 VSS VDD 16 480 20 VDD 532 VSS sky130_fd_sc_hd__dfstp_4 $T=91080 176800 0 0 $X=90890 $Y=176560
X3264 VSS VDD 416 497 20 VDD 285 VSS sky130_fd_sc_hd__dfstp_4 $T=92460 106080 0 0 $X=92270 $Y=105840
X3265 VSS VDD 17 496 20 VDD 510 VSS sky130_fd_sc_hd__dfstp_4 $T=93840 62560 0 0 $X=93650 $Y=62320
X3266 VSS VDD 17 523 20 VDD 525 VSS sky130_fd_sc_hd__dfstp_4 $T=99360 29920 0 0 $X=99170 $Y=29680
X3267 VSS VDD 17 725 20 VDD 719 VSS sky130_fd_sc_hd__dfstp_4 $T=135700 29920 1 0 $X=135510 $Y=26960
X3268 VSS VDD 16 601 20 VDD 801 VSS sky130_fd_sc_hd__dfstp_4 $T=149500 182240 0 0 $X=149310 $Y=182000
X3269 VSS VDD 16 660 20 VDD 823 VSS sky130_fd_sc_hd__dfstp_4 $T=152720 209440 0 0 $X=152530 $Y=209200
X3270 VSS VDD 17 792 20 VDD 872 VSS sky130_fd_sc_hd__dfstp_4 $T=158240 165920 0 0 $X=158050 $Y=165680
X3271 VSS VDD 16 563 20 VDD 855 VSS sky130_fd_sc_hd__dfstp_4 $T=158700 220320 0 0 $X=158510 $Y=220080
X3272 VSS VDD 17 809 20 VDD 887 VSS sky130_fd_sc_hd__dfstp_4 $T=161460 29920 1 0 $X=161270 $Y=26960
X3273 VSS VDD 17 833 20 VDD 945 VSS sky130_fd_sc_hd__dfstp_4 $T=176180 100640 0 0 $X=175990 $Y=100400
X3274 VSS VDD 17 854 20 VDD 947 VSS sky130_fd_sc_hd__dfstp_4 $T=176180 193120 0 0 $X=175990 $Y=192880
X3275 VSS VDD 17 847 20 VDD 956 VSS sky130_fd_sc_hd__dfstp_4 $T=179400 73440 0 0 $X=179210 $Y=73200
X3276 VSS VDD 17 880 20 VDD 969 VSS sky130_fd_sc_hd__dfstp_4 $T=183540 24480 0 0 $X=183350 $Y=24240
X3277 VSS VDD 315 271 331 347 316 328 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=58420 149600 1 0 $X=58230 $Y=146640
X3278 VSS VDD 575 605 585 531 594 461 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=110400 127840 1 0 $X=110210 $Y=124880
X3279 VSS VDD 640 635 675 685 686 424 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=126040 176800 0 0 $X=125850 $Y=176560
X3280 VSS VDD 718 712 346 728 734 233 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=136160 155040 1 0 $X=135970 $Y=152080
X3281 VSS VDD 736 726 716 710 742 652 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=138920 100640 1 0 $X=138730 $Y=97680
X3282 VSS VDD 902 519 887 930 884 890 VDD VSS sky130_fd_sc_hd__a32oi_4 $T=178940 40800 0 0 $X=178750 $Y=40560
X3283 VSS VDD 62 26 64 VDD 29 VSS sky130_fd_sc_hd__or3_4 $T=11960 95200 0 0 $X=11770 $Y=94960
X3284 VSS VDD 285 214 194 VDD 242 VSS sky130_fd_sc_hd__or3_4 $T=49680 100640 0 0 $X=49490 $Y=100400
X3285 VSS VDD 245 240 558 VDD 581 VSS sky130_fd_sc_hd__or3_4 $T=106720 209440 0 0 $X=106530 $Y=209200
X3286 VSS VDD 755 766 721 VDD 793 VSS sky130_fd_sc_hd__or3_4 $T=152260 138720 1 0 $X=152070 $Y=135760
X3287 VSS VDD 891 910 915 VDD 899 VSS sky130_fd_sc_hd__or3_4 $T=177100 144160 1 0 $X=176910 $Y=141200
X3288 VSS VDD 24 ICV_77 $T=8280 51680 0 0 $X=8090 $Y=51440
X3289 VSS VDD 66 ICV_77 $T=10580 106080 0 0 $X=10390 $Y=105840
X3290 VSS VDD 115 ICV_77 $T=20240 209440 0 0 $X=20050 $Y=209200
X3291 VSS VDD 94 ICV_77 $T=35880 127840 1 0 $X=35690 $Y=124880
X3292 VSS VDD 191 ICV_77 $T=61180 29920 1 0 $X=60990 $Y=26960
X3293 VSS VDD 3 ICV_77 $T=65320 84320 1 0 $X=65130 $Y=81360
X3294 VSS VDD 315 ICV_77 $T=77280 111520 1 0 $X=77090 $Y=108560
X3295 VSS VDD 429 ICV_77 $T=79580 165920 1 0 $X=79390 $Y=162960
X3296 VSS VDD 340 ICV_77 $T=84640 51680 1 0 $X=84450 $Y=48720
X3297 VSS VDD 583 ICV_77 $T=108560 225760 0 0 $X=108370 $Y=225520
X3298 VSS VDD 578 ICV_77 $T=149500 62560 0 0 $X=149310 $Y=62320
X3299 VSS VDD 778 ICV_77 $T=149500 187680 0 0 $X=149310 $Y=187440
X3300 VSS VDD 783 ICV_77 $T=160540 144160 0 0 $X=160350 $Y=143920
X3301 VSS VDD 788 ICV_77 $T=161460 51680 1 0 $X=161270 $Y=48720
X3302 VSS VDD 826 ICV_77 $T=161460 89760 1 0 $X=161270 $Y=86800
X3303 VSS VDD 891 ICV_77 $T=177100 138720 1 0 $X=176910 $Y=135760
X3304 VSS VDD 69 68 32 50 69 ICV_78 $T=9200 160480 1 0 $X=9010 $Y=157520
X3305 VSS VDD 504 518 SCAN_IN<11> 471 504 ICV_78 $T=93840 133280 1 0 $X=93650 $Y=130320
X3306 VSS VDD 529 606 529 574 559 ICV_78 $T=107640 68000 0 0 $X=107450 $Y=67760
X3307 VSS VDD 657 489 525 631 591 ICV_78 $T=119140 29920 0 0 $X=118950 $Y=29680
X3308 VSS VDD 671 692 671 290 647 ICV_78 $T=126500 214880 0 0 $X=126310 $Y=214640
X3309 VSS VDD 722 732 SCAN_IN<11> 661 711 ICV_78 $T=133400 116960 1 0 $X=133210 $Y=114000
X3310 VSS VDD 644 589 644 774 717 ICV_78 $T=148120 106080 0 0 $X=147930 $Y=105840
X3311 VSS VDD 920 904 878 418 853 ICV_78 $T=175260 19040 0 0 $X=175070 $Y=18800
X3312 VSS VDD 921 885 888 574 866 ICV_78 $T=175260 78880 0 0 $X=175070 $Y=78640
X3313 VSS VDD 915 910 846 891 894 ICV_78 $T=175260 138720 0 0 $X=175070 $Y=138480
X3314 VSS VDD 141 ICV_79 $T=25300 209440 1 0 $X=25110 $Y=206480
X3315 VSS VDD 185 ICV_79 $T=37260 46240 1 0 $X=37070 $Y=43280
X3316 VSS VDD 179 ICV_79 $T=45080 84320 0 0 $X=44890 $Y=84080
X3317 VSS VDD 301 ICV_79 $T=51520 214880 1 0 $X=51330 $Y=211920
X3318 VSS VDD 17 ICV_79 $T=93840 89760 0 0 $X=93650 $Y=89520
X3319 VSS VDD 638 ICV_79 $T=120060 68000 1 0 $X=119870 $Y=65040
X3320 VSS VDD 795 ICV_79 $T=161460 198560 1 0 $X=161270 $Y=195600
X3321 VSS VDD 846 ICV_79 $T=165140 133280 0 0 $X=164950 $Y=133040
X3322 VSS VDD 418 ICV_79 $T=174340 24480 1 0 $X=174150 $Y=21520
X3323 VSS VDD ICV_80 $T=17480 225760 1 0 $X=17290 $Y=222800
X3324 VSS VDD ICV_80 $T=31280 106080 0 0 $X=31090 $Y=105840
X3325 VSS VDD ICV_80 $T=59340 35360 0 0 $X=59150 $Y=35120
X3326 VSS VDD ICV_80 $T=59340 62560 0 0 $X=59150 $Y=62320
X3327 VSS VDD ICV_80 $T=59340 133280 0 0 $X=59150 $Y=133040
X3328 VSS VDD ICV_80 $T=73600 214880 1 0 $X=73410 $Y=211920
X3329 VSS VDD ICV_80 $T=87400 46240 0 0 $X=87210 $Y=46000
X3330 VSS VDD ICV_80 $T=87400 68000 0 0 $X=87210 $Y=67760
X3331 VSS VDD ICV_80 $T=101660 46240 1 0 $X=101470 $Y=43280
X3332 VSS VDD ICV_80 $T=143520 116960 0 0 $X=143330 $Y=116720
X3333 VSS VDD ICV_80 $T=174340 13600 1 0 $X=174150 $Y=10640
X3334 VSS VDD 328 319 335 329 336 VDD 200 VSS sky130_fd_sc_hd__o41a_4 $T=62100 160480 1 0 $X=61910 $Y=157520
X3335 VSS VDD 890 906 874 869 897 VDD 707 VSS sky130_fd_sc_hd__o41a_4 $T=172960 40800 1 0 $X=172770 $Y=37840
X3336 VSS VDD 287 294 303 322 VDD 107 VSS sky130_fd_sc_hd__nor4_4 $T=50600 40800 1 0 $X=50410 $Y=37840
X3337 VSS VDD 366 375 362 107 VDD 3 VSS sky130_fd_sc_hd__nor4_4 $T=64400 68000 0 0 $X=64210 $Y=67760
X3338 VSS VDD 114 230 404 409 VDD 437 VSS sky130_fd_sc_hd__nor4_4 $T=77280 144160 1 0 $X=77090 $Y=141200
X3339 VSS VDD 458 617 561 109 VDD 662 VSS sky130_fd_sc_hd__nor4_4 $T=118680 149600 1 0 $X=118490 $Y=146640
X3340 VSS VDD 458 625 610 109 VDD 667 VSS sky130_fd_sc_hd__nor4_4 $T=119140 155040 0 0 $X=118950 $Y=154800
X3341 VSS VDD 607 672 860 898 VDD 891 VSS sky130_fd_sc_hd__nor4_4 $T=171120 106080 1 0 $X=170930 $Y=103120
X3342 VSS VDD 120 ICV_81 $T=30820 111520 0 0 $X=30630 $Y=111280
X3343 VSS VDD 275 ICV_81 $T=58880 68000 0 0 $X=58690 $Y=67760
X3344 VSS VDD 315 ICV_81 $T=58880 122400 0 0 $X=58690 $Y=122160
X3345 VSS VDD 489 ICV_81 $T=115000 40800 0 0 $X=114810 $Y=40560
X3346 VSS VDD 573 ICV_81 $T=115000 84320 0 0 $X=114810 $Y=84080
X3347 VSS VDD 321 ICV_81 $T=115000 187680 0 0 $X=114810 $Y=187440
X3348 VSS VDD 865 ICV_81 $T=171120 24480 0 0 $X=170930 $Y=24240
X3349 VSS VDD 607 ICV_81 $T=171120 100640 0 0 $X=170930 $Y=100400
X3350 VSS VDD 102 ICV_82 $T=16560 133280 1 0 $X=16370 $Y=130320
X3351 VSS VDD 194 ICV_82 $T=30360 100640 0 0 $X=30170 $Y=100400
X3352 VSS VDD 87 ICV_82 $T=30360 193120 0 0 $X=30170 $Y=192880
X3353 VSS VDD 197 ICV_82 $T=30360 209440 0 0 $X=30170 $Y=209200
X3354 VSS VDD 269 ICV_82 $T=44620 171360 1 0 $X=44430 $Y=168400
X3355 VSS VDD 121 ICV_82 $T=86480 35360 0 0 $X=86290 $Y=35120
X3356 VSS VDD 184 ICV_82 $T=114540 214880 0 0 $X=114350 $Y=214640
X3357 VSS VDD 894 ICV_82 $T=170660 144160 0 0 $X=170470 $Y=143920
X3358 VSS VDD 11 29 28 VDD 45 VSS sky130_fd_sc_hd__and3_4 $T=7820 100640 0 0 $X=7630 $Y=100400
X3359 VSS VDD 11 27 66 VDD 56 VSS sky130_fd_sc_hd__and3_4 $T=10580 106080 1 0 $X=10390 $Y=103120
X3360 VSS VDD 11 44 36 VDD 86 VSS sky130_fd_sc_hd__and3_4 $T=11040 95200 1 0 $X=10850 $Y=92240
X3361 VSS VDD 11 74 63 VDD 89 VSS sky130_fd_sc_hd__and3_4 $T=11500 78880 1 0 $X=11310 $Y=75920
X3362 VSS VDD 102 96 104 VDD 76 VSS sky130_fd_sc_hd__and3_4 $T=18860 176800 0 0 $X=18670 $Y=176560
X3363 VSS VDD 565 584 577 VDD 542 VSS sky130_fd_sc_hd__and3_4 $T=108100 73440 0 0 $X=107910 $Y=73200
X3364 VSS VDD 747 SCAN_IN<0> 863 VDD 901 VSS sky130_fd_sc_hd__and3_4 $T=170200 220320 1 0 $X=170010 $Y=217360
X3365 VSS VDD 20 169 212 ICV_83 $T=55660 13600 0 0 $X=55470 $Y=13360
X3366 VSS VDD 339 378 349 ICV_83 $T=69920 182240 1 0 $X=69730 $Y=179280
X3367 VSS VDD 58 451 401 ICV_83 $T=83720 193120 0 0 $X=83530 $Y=192880
X3368 VSS VDD 502 501 510 ICV_83 $T=97980 57120 1 0 $X=97790 $Y=54160
X3369 VSS VDD 509 SCAN_IN<21> 565 ICV_83 $T=106720 84320 0 0 $X=106530 $Y=84080
X3370 VSS VDD 603 573 570 ICV_83 $T=111780 24480 0 0 $X=111590 $Y=24240
X3371 VSS VDD 579 301 92 ICV_83 $T=111780 209440 0 0 $X=111590 $Y=209200
X3372 VSS VDD 611 612 623 ICV_83 $T=114540 24480 1 0 $X=114350 $Y=21520
X3373 VSS VDD 640 675 686 ICV_83 $T=126040 176800 1 0 $X=125850 $Y=173840
X3374 VSS VDD 867 861 848 ICV_83 $T=167900 89760 0 0 $X=167710 $Y=89520
X3375 VSS VDD 868 877 558 ICV_83 $T=167900 209440 0 0 $X=167710 $Y=209200
X3376 VSS VDD 78 83 40 76 92 51 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=11960 187680 0 0 $X=11770 $Y=187440
X3377 VSS VDD 126 123 97 111 92 52 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=21160 204000 1 0 $X=20970 $Y=201040
X3378 VSS VDD 314 291 320 313 321 311 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=54280 204000 1 0 $X=54090 $Y=201040
X3379 VSS VDD 384 367 381 380 346 352 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=69000 106080 0 0 $X=68810 $Y=105840
X3380 VSS VDD 459 457 446 469 321 480 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=86020 193120 1 0 $X=85830 $Y=190160
X3381 VSS VDD 463 483 477 447 401 495 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=88780 220320 1 0 $X=88590 $Y=217360
X3382 VSS VDD 524 527 559 542 551 496 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=105340 73440 1 0 $X=105150 $Y=70480
X3383 VSS VDD 543 546 540 539 321 601 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=106720 193120 1 0 $X=106530 $Y=190160
X3384 VSS VDD 564 571 593 587 551 523 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=107180 40800 1 0 $X=106990 $Y=37840
X3385 VSS VDD 602 621 627 626 321 660 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=119140 204000 0 0 $X=118950 $Y=203760
X3386 VSS VDD 782 781 797 805 698 809 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=153180 40800 0 0 $X=152990 $Y=40560
X3387 VSS VDD 811 806 812 832 698 833 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=161460 100640 1 0 $X=161270 $Y=97680
X3388 VSS VDD 814 828 852 839 787 871 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=163760 155040 1 0 $X=163570 $Y=152080
X3389 VSS VDD 825 831 866 850 698 847 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=164220 78880 1 0 $X=164030 $Y=75920
X3390 VSS VDD 827 858 849 856 698 854 VDD VSS sky130_fd_sc_hd__o32ai_4 $T=164680 116960 1 0 $X=164490 $Y=114000
X3391 VSS VDD 63 11 74 ICV_84 $T=12880 73440 0 0 $X=12690 $Y=73200
X3392 VSS VDD 167 19 133 ICV_84 $T=23920 29920 1 0 $X=23730 $Y=26960
X3393 VSS VDD 92 126 87 ICV_84 $T=24840 198560 0 0 $X=24650 $Y=198320
X3394 VSS VDD 94 20 293 ICV_84 $T=49220 171360 0 0 $X=49030 $Y=171120
X3395 VSS VDD 132 286 271 ICV_84 $T=49220 176800 0 0 $X=49030 $Y=176560
X3396 VSS VDD 416 20 434 ICV_84 $T=78200 35360 0 0 $X=78010 $Y=35120
X3397 VSS VDD 494 230 449 ICV_84 $T=94300 138720 1 0 $X=94110 $Y=135760
X3398 VSS VDD 456 20 569 ICV_84 $T=104420 155040 0 0 $X=104230 $Y=154800
X3399 VSS VDD 466 346 592 ICV_84 $T=108100 111520 0 0 $X=107910 $Y=111280
X3400 VSS VDD 456 20 709 ICV_84 $T=132480 73440 0 0 $X=132290 $Y=73200
X3401 VSS VDD 745 731 453 ICV_84 $T=137540 62560 0 0 $X=137350 $Y=62320
X3402 VSS VDD 537 633 786 ICV_84 $T=148580 193120 0 0 $X=148390 $Y=192880
X3403 VSS VDD 703 830 730 ICV_84 $T=164220 40800 0 0 $X=164030 $Y=40560
X3404 VSS VDD 843 845 838 ICV_84 $T=164680 62560 0 0 $X=164490 $Y=62320
X3405 VSS VDD 59 65 48 48 ICV_85 $T=6900 193120 1 0 $X=6710 $Y=190160
X3406 VSS VDD 191 124 209 154 ICV_85 $T=33580 19040 1 0 $X=33390 $Y=16080
X3407 VSS VDD 55 276 392 55 ICV_85 $T=69460 73440 0 0 $X=69270 $Y=73200
X3408 VSS VDD 370 7 381 370 ICV_85 $T=75440 100640 0 0 $X=75250 $Y=100400
X3409 VSS VDD 400 418 425 SCAN_IN<7> ICV_85 $T=75440 149600 0 0 $X=75250 $Y=149360
X3410 VSS VDD SCAN_IN<13> 680 485 680 ICV_85 $T=134320 144160 0 0 $X=134130 $Y=143920
X3411 VSS VDD 727 SCAN_IN<12> 739 727 ICV_85 $T=135240 138720 0 0 $X=135050 $Y=138480
X3412 VSS VDD 788 796 780 788 ICV_85 $T=154100 29920 0 0 $X=153910 $Y=29680
X3413 VSS VDD 769 790 828 787 ICV_85 $T=161920 149600 0 0 $X=161730 $Y=149360
X3414 VSS VDD 848 574 812 848 ICV_85 $T=163300 95200 0 0 $X=163110 $Y=94960
X3415 VSS VDD 64 62 64 27 ICV_86 $T=19780 95200 0 0 $X=19590 $Y=94960
X3416 VSS VDD 119 81 119 85 ICV_86 $T=22080 57120 0 0 $X=21890 $Y=56880
X3417 VSS VDD 168 85 61 157 ICV_86 $T=23460 46240 1 0 $X=23270 $Y=43280
X3418 VSS VDD 154 107 154 108 ICV_86 $T=24840 62560 0 0 $X=24650 $Y=62320
X3419 VSS VDD 330 284 275 289 ICV_86 $T=54740 68000 1 0 $X=54550 $Y=65040
X3420 VSS VDD 331 353 331 286 ICV_86 $T=64860 176800 0 0 $X=64670 $Y=176560
X3421 VSS VDD 506 491 506 470 ICV_86 $T=94760 198560 0 0 $X=94570 $Y=198320
X3422 VSS VDD 512 512 506 482 ICV_86 $T=97060 171360 1 0 $X=96870 $Y=168400
X3423 VSS VDD 506 476 506 600 ICV_86 $T=109020 165920 0 0 $X=108830 $Y=165680
X3424 VSS VDD SCAN_IN<20> SCAN_IN<20> 598 588 ICV_86 $T=110860 100640 0 0 $X=110670 $Y=100400
X3425 VSS VDD 671 708 671 692 ICV_86 $T=136620 225760 1 0 $X=136430 $Y=222800
X3426 VSS VDD 622 578 622 744 ICV_86 $T=138920 57120 0 0 $X=138730 $Y=56880
X3427 VSS VDD 521 824 521 843 ICV_86 $T=161920 62560 1 0 $X=161730 $Y=59600
X3428 VSS VDD 75 131 118 VDD 103 VSS sky130_fd_sc_hd__a21boi_4 $T=21160 165920 1 0 $X=20970 $Y=162960
X3429 VSS VDD 133 117 128 VDD 134 VSS sky130_fd_sc_hd__a21boi_4 $T=23000 35360 1 0 $X=22810 $Y=32400
X3430 VSS VDD 146 151 145 VDD 162 VSS sky130_fd_sc_hd__a21boi_4 $T=24380 220320 1 0 $X=24190 $Y=217360
X3431 VSS VDD 267 242 266 VDD 229 VSS sky130_fd_sc_hd__a21boi_4 $T=47380 89760 0 0 $X=47190 $Y=89520
X3432 VSS VDD 297 343 349 VDD 359 VSS sky130_fd_sc_hd__a21boi_4 $T=63020 220320 0 0 $X=62830 $Y=220080
X3433 VSS VDD 612 655 623 VDD 611 VSS sky130_fd_sc_hd__a21boi_4 $T=119140 19040 0 0 $X=118950 $Y=18800
X3434 VSS VDD 684 694 608 VDD 714 VSS sky130_fd_sc_hd__a21boi_4 $T=132940 35360 0 0 $X=132750 $Y=35120
X3435 VSS VDD 796 802 810 VDD 824 VSS sky130_fd_sc_hd__a21boi_4 $T=160080 57120 0 0 $X=159890 $Y=56880
X3436 VSS VDD 13 VDD 31 VSS sky130_fd_sc_hd__clkbuf_16 $T=7820 138720 1 0 $X=7630 $Y=135760
X3437 VSS VDD 60 VDD 171 VSS sky130_fd_sc_hd__clkbuf_16 $T=39100 68000 0 0 $X=38910 $Y=67760
X3438 VSS VDD 277 VDD 216 VSS sky130_fd_sc_hd__clkbuf_16 $T=49680 73440 0 0 $X=49490 $Y=73200
X3439 VSS VDD 299 VDD 94 VSS sky130_fd_sc_hd__clkbuf_16 $T=51980 133280 1 0 $X=51790 $Y=130320
X3440 VSS VDD 135 VDD 299 VSS sky130_fd_sc_hd__clkbuf_16 $T=77280 127840 1 0 $X=77090 $Y=124880
X3441 VSS VDD CLK_IN VDD 277 VSS sky130_fd_sc_hd__clkbuf_16 $T=91080 13600 0 0 $X=90890 $Y=13360
X3442 VSS VDD 299 VDD 456 VSS sky130_fd_sc_hd__clkbuf_16 $T=91080 116960 0 0 $X=90890 $Y=116720
X3443 VSS VDD 614 VDD 416 VSS sky130_fd_sc_hd__clkbuf_16 $T=116840 78880 1 0 $X=116650 $Y=75920
X3444 VSS VDD 487 VDD 614 VSS sky130_fd_sc_hd__clkbuf_16 $T=142600 84320 1 0 $X=142410 $Y=81360
X3445 VSS VDD 614 VDD 844 VSS sky130_fd_sc_hd__clkbuf_16 $T=155940 78880 0 0 $X=155750 $Y=78640
X3446 VSS VDD 158 114 137 ICV_87 $T=24380 133280 0 0 $X=24190 $Y=133040
X3447 VSS VDD 94 20 306 ICV_87 $T=53820 116960 0 0 $X=53630 $Y=116720
X3448 VSS VDD 220 342 344 ICV_87 $T=61640 62560 1 0 $X=61450 $Y=59600
X3449 VSS VDD 360 354 369 ICV_87 $T=66700 78880 1 0 $X=66510 $Y=75920
X3450 VSS VDD 416 20 435 ICV_87 $T=78660 57120 0 0 $X=78470 $Y=56880
X3451 VSS VDD 416 20 445 ICV_87 $T=81880 40800 0 0 $X=81690 $Y=40560
X3452 VSS VDD 568 561 471 ICV_87 $T=109940 149600 0 0 $X=109750 $Y=149360
X3453 VSS VDD 800 793 794 ICV_87 $T=152720 160480 1 0 $X=152530 $Y=157520
X3454 VSS VDD 683 20 20 ICV_87 $T=152720 214880 1 0 $X=152530 $Y=211920
X3455 VSS VDD ICV_88 $T=34040 149600 1 0 $X=33850 $Y=146640
X3456 VSS VDD ICV_88 $T=77280 13600 1 0 $X=77090 $Y=10640
X3457 VSS VDD ICV_89 $T=20240 225760 0 0 $X=20050 $Y=225520
X3458 VSS VDD ICV_89 $T=48760 13600 1 0 $X=48570 $Y=10640
X3459 VSS VDD ICV_89 $T=48760 225760 0 0 $X=48570 $Y=225520
X3460 VSS VDD ICV_89 $T=120060 225760 0 0 $X=119870 $Y=225520
X3461 VSS VDD ICV_89 $T=148580 225760 0 0 $X=148390 $Y=225520
X3462 VSS VDD 284 267 276 VDD 181 VSS sky130_fd_sc_hd__a21bo_4 $T=49220 78880 1 0 $X=49030 $Y=75920
X3463 VSS VDD 289 284 275 VDD 193 VSS sky130_fd_sc_hd__a21bo_4 $T=49680 62560 0 0 $X=49490 $Y=62320
X3464 VSS VDD 379 289 330 VDD 351 VSS sky130_fd_sc_hd__a21bo_4 $T=69000 57120 0 0 $X=68810 $Y=56880
X3465 VSS VDD 391 379 373 VDD 350 VSS sky130_fd_sc_hd__a21bo_4 $T=77280 51680 1 0 $X=77090 $Y=48720
X3466 VSS VDD 762 764 628 VDD 655 VSS sky130_fd_sc_hd__a21bo_4 $T=147660 19040 1 0 $X=147470 $Y=16080
X3467 VSS VDD 49 70 VDD 35 VSS sky130_fd_sc_hd__xor2_4 $T=9200 13600 0 0 $X=9010 $Y=13360
X3468 VSS VDD 67 82 VDD 90 VSS sky130_fd_sc_hd__xor2_4 $T=10580 149600 0 0 $X=10390 $Y=149360
X3469 VSS VDD 252 292 VDD 256 VSS sky130_fd_sc_hd__xor2_4 $T=49220 160480 1 0 $X=49030 $Y=157520
X3470 VSS VDD 508 514 VDD 570 VSS sky130_fd_sc_hd__xor2_4 $T=97520 24480 0 0 $X=97330 $Y=24240
X3471 VSS VDD 697 724 VDD 764 VSS sky130_fd_sc_hd__xor2_4 $T=147660 13600 0 0 $X=147470 $Y=13360
X3472 VSS VDD 485 494 504 449 230 VDD 488 VSS sky130_fd_sc_hd__a2111o_4 $T=92460 133280 0 0 $X=92270 $Y=133040
X3473 VSS VDD 237 665 653 641 620 VDD 645 VSS sky130_fd_sc_hd__a2111o_4 $T=124200 187680 0 0 $X=124010 $Y=187440
X3474 VSS VDD 702 711 717 672 449 VDD 729 VSS sky130_fd_sc_hd__a2111o_4 $T=133400 111520 1 0 $X=133210 $Y=108560
X3475 VSS VDD 472 517 518 436 VDD 498 VSS sky130_fd_sc_hd__nand4_4 $T=95220 127840 0 0 $X=95030 $Y=127600
X3476 VSS VDD 704 648 710 664 VDD 720 VSS sky130_fd_sc_hd__nand4_4 $T=133400 106080 1 0 $X=133210 $Y=103120
X3477 VSS VDD 38 VDD 13 VSS sky130_fd_sc_hd__clkbuf_4 $T=8280 133280 1 0 $X=8090 $Y=130320
X3478 VSS VDD 38 VDD 60 VSS sky130_fd_sc_hd__clkbuf_4 $T=8740 19040 1 0 $X=8550 $Y=16080
X3479 VSS VDD 121 VDD 135 VSS sky130_fd_sc_hd__clkbuf_4 $T=21160 122400 0 0 $X=20970 $Y=122160
X3480 VSS VDD 121 VDD 487 VSS sky130_fd_sc_hd__clkbuf_4 $T=91080 35360 0 0 $X=90890 $Y=35120
X3481 VSS VDD 31 12 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=7820 127840 1 0 $X=7630 $Y=124880
X3482 VSS VDD 31 14 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=7820 149600 0 0 $X=7630 $Y=149360
X3483 VSS VDD 171 10 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=29440 68000 0 0 $X=29250 $Y=67760
X3484 VSS VDD 216 38 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=36800 73440 0 0 $X=36610 $Y=73200
X3485 VSS VDD 171 212 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=45080 73440 1 0 $X=44890 $Y=70480
X3486 VSS VDD 216 121 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=57040 78880 0 0 $X=56850 $Y=78640
X3487 18 VDD VSS sky130_fd_sc_hd__conb_1 $T=7820 220320 1 0 $X=7630 $Y=217360
X3488 41 VDD VSS sky130_fd_sc_hd__conb_1 $T=8740 225760 1 0 $X=8550 $Y=222800
X3489 VSS VDD ICV_90 $T=5520 13600 1 0 $X=5330 $Y=10640
X3490 VSS VDD ICV_90 $T=5520 13600 0 0 $X=5330 $Y=13360
X3491 VSS VDD ICV_90 $T=5520 19040 1 0 $X=5330 $Y=16080
X3492 VSS VDD ICV_90 $T=5520 68000 0 0 $X=5330 $Y=67760
X3493 VSS VDD ICV_90 $T=5520 160480 1 0 $X=5330 $Y=157520
X3494 VSS VDD ICV_90 $T=5520 165920 1 0 $X=5330 $Y=162960
X3495 VSS VDD ICV_90 $T=5520 165920 0 0 $X=5330 $Y=165680
X3496 VSS VDD ICV_90 $T=5520 193120 0 0 $X=5330 $Y=192880
X3497 VSS VDD ICV_90 $T=5520 220320 0 0 $X=5330 $Y=220080
X3498 VSS VDD ICV_90 $T=5520 225760 1 0 $X=5330 $Y=222800
.ENDS
***************************************
