* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_6000626648221
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_CDNS_6000626648219 2 3 4
** N=24 EP=3 IP=6 FDC=1
*.SEEDPROM
M0 4 3 2 2 pshort L=0.15 W=7 m=1 r=46.6667 a=1.05 p=14.3 mult=1 $X=0 $Y=0 $D=79
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_6000626648224
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_CDNS_6000626648222 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 4 2 3 1 nshort L=0.15 W=7 m=1 r=46.6667 a=1.05 p=14.3 mult=1 $X=0 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT NAND GND INP1 INP2 VDD OUT
** N=44 EP=5 IP=16 FDC=6
X0 GND VDD Dpar a=12.6592 p=18.16 m=1 $[nwdiode] $X=2130 $Y=9720 $D=191
X1 GND VDD Dpar a=12.6592 p=18.16 m=1 $[nwdiode] $X=5305 $Y=9705 $D=191
X2 VDD INP1 OUT pfet_CDNS_6000626648219 $T=3255 9900 0 0 $X=2130 $Y=9720
X3 VDD INP2 OUT pfet_CDNS_6000626648219 $T=6430 9885 0 0 $X=5305 $Y=9705
X4 GND INP1 6 OUT nfet_CDNS_6000626648222 $T=3255 1885 0 0 $X=2865 $Y=1755
X5 GND INP2 GND 6 nfet_CDNS_6000626648222 $T=6580 1885 1 180 $X=6040 $Y=1755
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_600062664826
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_600062664822
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_600062664827
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT Inverter0 GND VDD INP OUT
** N=32 EP=4 IP=11 FDC=4
M0 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3140 $Y=1490 $D=9
M1 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2915 $Y=7755 $D=79
M2 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3345 $Y=7755 $D=79
X3 GND VDD Dpar a=11.524 p=15.02 m=1 $[nwdiode] $X=1790 $Y=7575 $D=191
.ENDS
***************************************
.SUBCKT ICV_1
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_600062664823
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT Inverter2 GND VDD INP OUT
** N=32 EP=4 IP=31 FDC=28
M0 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2210 $Y=1130 $D=9
M1 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2640 $Y=1130 $D=9
M2 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3070 $Y=1130 $D=9
M3 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3500 $Y=1130 $D=9
M4 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3930 $Y=1130 $D=9
M5 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4360 $Y=1130 $D=9
M6 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4790 $Y=1130 $D=9
M7 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5220 $Y=1130 $D=9
M8 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5650 $Y=1130 $D=9
M9 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1985 $Y=7395 $D=79
M10 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2415 $Y=7395 $D=79
M11 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2845 $Y=7395 $D=79
M12 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3275 $Y=7395 $D=79
M13 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3705 $Y=7395 $D=79
M14 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4135 $Y=7395 $D=79
M15 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4565 $Y=7395 $D=79
M16 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4995 $Y=7395 $D=79
M17 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5425 $Y=7395 $D=79
M18 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5855 $Y=7395 $D=79
M19 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6285 $Y=7395 $D=79
M20 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6715 $Y=7395 $D=79
M21 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7145 $Y=7395 $D=79
M22 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7575 $Y=7395 $D=79
M23 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8005 $Y=7395 $D=79
M24 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8435 $Y=7395 $D=79
M25 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8865 $Y=7395 $D=79
M26 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=9295 $Y=7395 $D=79
X27 GND VDD Dpar a=48.4008 p=28.78 m=1 $[nwdiode] $X=860 $Y=7215 $D=191
.ENDS
***************************************
.SUBCKT pfet_CDNS_600062664828 2 3 4
** N=7 EP=3 IP=0 FDC=1
*.SEEDPROM
M0 3 3 4 2 pshort L=8 W=0.55 m=1 r=0.06875 a=4.4 p=17.1 mult=1 $X=0 $Y=0 $D=79
.ENDS
***************************************
.SUBCKT Receiver GND VDD INP CLK OUT_B OUT
** N=47 EP=6 IP=81 FDC=98
M0 5 INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5690 $Y=12530 $D=9
M1 GND INP 5 GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6120 $Y=12530 $D=9
M2 5 INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6550 $Y=12530 $D=9
M3 5 INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5465 $Y=18795 $D=79
M4 VDD INP 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5895 $Y=18795 $D=79
M5 5 INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6325 $Y=18795 $D=79
M6 VDD INP 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6755 $Y=18795 $D=79
M7 5 INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7185 $Y=18795 $D=79
M8 VDD INP 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7615 $Y=18795 $D=79
X9 GND VDD Dpar a=8.7087 p=20.96 m=1 $[nwdiode] $X=1885 $Y=18755 $D=191
X10 GND VDD Dpar a=20.7432 p=18.46 m=1 $[nwdiode] $X=4340 $Y=18615 $D=191
X11 GND VDD Dpar a=8.7087 p=20.96 m=1 $[nwdiode] $X=9500 $Y=18810 $D=191
X12 GND 6 CLK VDD 15 NAND $T=25500 17975 0 0 $X=26890 $Y=18460
X13 GND 7 CLK VDD 14 NAND $T=25505 -25 0 0 $X=26895 $Y=460
X14 GND 14 10 VDD 9 NAND $T=33045 120 0 0 $X=34435 $Y=605
X15 GND 15 9 VDD 10 NAND $T=33155 18005 0 0 $X=34545 $Y=18490
X16 GND 9 11 VDD 16 NAND $T=41280 120 0 0 $X=42670 $Y=605
X17 GND 10 11 VDD 17 NAND $T=41390 18005 0 0 $X=42780 $Y=18490
X18 GND 16 OUT VDD OUT_B NAND $T=52015 120 0 0 $X=53405 $Y=605
X19 GND 17 OUT_B VDD OUT NAND $T=52125 18005 0 0 $X=53515 $Y=18490
X25 GND VDD 6 7 Inverter0 $T=21660 11035 0 0 $X=22845 $Y=11745
X26 GND VDD CLK 11 Inverter0 $T=47900 11035 0 0 $X=49085 $Y=11745
X31 GND VDD 5 6 Inverter2 $T=11225 11395 0 0 $X=11480 $Y=11745
X32 VDD 3 INP pfet_CDNS_600062664828 $T=2615 19880 0 90 $X=1885 $Y=18755
X33 VDD 5 3 pfet_CDNS_600062664828 $T=9680 27255 0 270 $X=9500 $Y=18810
.ENDS
***************************************
