* NGSPICE file created from serializer_unit_cell_1.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

.subckt serializer_unit_cell_1 CLK COMPLETE COUNT[0] COUNT[1] COUNT[2] COUNT[3] COUNT[4]
+ COUNT[5] INTERNAL_FINISH PAR_IN1[0] PAR_IN1[10] PAR_IN1[11] PAR_IN1[12] PAR_IN1[13]
+ PAR_IN1[14] PAR_IN1[15] PAR_IN1[16] PAR_IN1[17] PAR_IN1[18] PAR_IN1[19] PAR_IN1[1]
+ PAR_IN1[20] PAR_IN1[21] PAR_IN1[22] PAR_IN1[23] PAR_IN1[24] PAR_IN1[25] PAR_IN1[26]
+ PAR_IN1[27] PAR_IN1[28] PAR_IN1[29] PAR_IN1[2] PAR_IN1[30] PAR_IN1[31] PAR_IN1[3]
+ PAR_IN1[4] PAR_IN1[5] PAR_IN1[6] PAR_IN1[7] PAR_IN1[8] PAR_IN1[9] PAR_IN2[0] PAR_IN2[10]
+ PAR_IN2[11] PAR_IN2[12] PAR_IN2[13] PAR_IN2[14] PAR_IN2[15] PAR_IN2[16] PAR_IN2[17]
+ PAR_IN2[18] PAR_IN2[19] PAR_IN2[1] PAR_IN2[20] PAR_IN2[21] PAR_IN2[22] PAR_IN2[23]
+ PAR_IN2[24] PAR_IN2[25] PAR_IN2[26] PAR_IN2[27] PAR_IN2[28] PAR_IN2[29] PAR_IN2[2]
+ PAR_IN2[30] PAR_IN2[31] PAR_IN2[3] PAR_IN2[4] PAR_IN2[5] PAR_IN2[6] PAR_IN2[7] PAR_IN2[8]
+ PAR_IN2[9] PAR_IN3[0] PAR_IN3[10] PAR_IN3[11] PAR_IN3[12] PAR_IN3[13] PAR_IN3[14]
+ PAR_IN3[15] PAR_IN3[16] PAR_IN3[17] PAR_IN3[18] PAR_IN3[19] PAR_IN3[1] PAR_IN3[20]
+ PAR_IN3[21] PAR_IN3[22] PAR_IN3[23] PAR_IN3[24] PAR_IN3[25] PAR_IN3[26] PAR_IN3[27]
+ PAR_IN3[28] PAR_IN3[29] PAR_IN3[2] PAR_IN3[30] PAR_IN3[31] PAR_IN3[3] PAR_IN3[4]
+ PAR_IN3[5] PAR_IN3[6] PAR_IN3[7] PAR_IN3[8] PAR_IN3[9] PAR_IN4[0] PAR_IN4[10] PAR_IN4[11]
+ PAR_IN4[12] PAR_IN4[13] PAR_IN4[14] PAR_IN4[15] PAR_IN4[16] PAR_IN4[17] PAR_IN4[18]
+ PAR_IN4[19] PAR_IN4[1] PAR_IN4[20] PAR_IN4[21] PAR_IN4[22] PAR_IN4[23] PAR_IN4[24]
+ PAR_IN4[25] PAR_IN4[26] PAR_IN4[27] PAR_IN4[28] PAR_IN4[29] PAR_IN4[2] PAR_IN4[30]
+ PAR_IN4[31] PAR_IN4[3] PAR_IN4[4] PAR_IN4[5] PAR_IN4[6] PAR_IN4[7] PAR_IN4[8] PAR_IN4[9]
+ PAR_IN5[0] PAR_IN5[10] PAR_IN5[11] PAR_IN5[12] PAR_IN5[13] PAR_IN5[14] PAR_IN5[15]
+ PAR_IN5[16] PAR_IN5[17] PAR_IN5[18] PAR_IN5[19] PAR_IN5[1] PAR_IN5[20] PAR_IN5[21]
+ PAR_IN5[22] PAR_IN5[23] PAR_IN5[24] PAR_IN5[25] PAR_IN5[26] PAR_IN5[27] PAR_IN5[28]
+ PAR_IN5[29] PAR_IN5[2] PAR_IN5[30] PAR_IN5[31] PAR_IN5[3] PAR_IN5[4] PAR_IN5[5]
+ PAR_IN5[6] PAR_IN5[7] PAR_IN5[8] PAR_IN5[9] PAR_IN6[0] PAR_IN6[10] PAR_IN6[11] PAR_IN6[12]
+ PAR_IN6[13] PAR_IN6[14] PAR_IN6[15] PAR_IN6[16] PAR_IN6[17] PAR_IN6[18] PAR_IN6[19]
+ PAR_IN6[1] PAR_IN6[20] PAR_IN6[21] PAR_IN6[22] PAR_IN6[23] PAR_IN6[24] PAR_IN6[25]
+ PAR_IN6[26] PAR_IN6[27] PAR_IN6[28] PAR_IN6[29] PAR_IN6[2] PAR_IN6[30] PAR_IN6[31]
+ PAR_IN6[3] PAR_IN6[4] PAR_IN6[5] PAR_IN6[6] PAR_IN6[7] PAR_IN6[8] PAR_IN6[9] PAR_IN7[0]
+ PAR_IN7[10] PAR_IN7[11] PAR_IN7[12] PAR_IN7[13] PAR_IN7[14] PAR_IN7[15] PAR_IN7[16]
+ PAR_IN7[17] PAR_IN7[18] PAR_IN7[19] PAR_IN7[1] PAR_IN7[20] PAR_IN7[21] PAR_IN7[22]
+ PAR_IN7[23] PAR_IN7[24] PAR_IN7[25] PAR_IN7[26] PAR_IN7[27] PAR_IN7[28] PAR_IN7[29]
+ PAR_IN7[2] PAR_IN7[30] PAR_IN7[31] PAR_IN7[3] PAR_IN7[4] PAR_IN7[5] PAR_IN7[6] PAR_IN7[7]
+ PAR_IN7[8] PAR_IN7[9] PAR_IN8[0] PAR_IN8[10] PAR_IN8[11] PAR_IN8[12] PAR_IN8[13]
+ PAR_IN8[14] PAR_IN8[15] PAR_IN8[16] PAR_IN8[17] PAR_IN8[18] PAR_IN8[19] PAR_IN8[1]
+ PAR_IN8[20] PAR_IN8[21] PAR_IN8[22] PAR_IN8[23] PAR_IN8[24] PAR_IN8[25] PAR_IN8[26]
+ PAR_IN8[27] PAR_IN8[28] PAR_IN8[29] PAR_IN8[2] PAR_IN8[30] PAR_IN8[31] PAR_IN8[3]
+ PAR_IN8[4] PAR_IN8[5] PAR_IN8[6] PAR_IN8[7] PAR_IN8[8] PAR_IN8[9] READY RESET SAMPLE_COUNT[0]
+ SAMPLE_COUNT[1] SAMPLE_COUNT[2] SAMPLE_COUNT[3] SERIAL_OUT VDD VSS
XFILLER_39_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_19 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_317 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0717__B1 _0643_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_280 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0613__A _0842_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_188 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0986__C _0985_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0708__B1 _0707_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_45 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0947__B1 _0946_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0985_ _0985_/A _0985_/B _0982_/X _0984_/X _0985_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0523__A _0522_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_29 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_214 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_10_169 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0938__B1 _0937_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_65 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_53_94 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_250 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_280 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0608__A _0608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0929__B1 _0792_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0770_ PAR_IN6[29] _0597_/X _0770_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0641__A2 _0606_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0997__B _0988_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_195 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0518__A _0518_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_239 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_291 VSS VDD sky130_fd_sc_hd__fill_2
X_0968_ PAR_IN2[28] _0925_/B _0968_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0899_ _0510_/X _0899_/B _0898_/X _0900_/C VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_23_250 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_206 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_217 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_228 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0871__A2 _0646_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0610__B _0610_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_176 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_143 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_250 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_294 VSS VDD sky130_fd_sc_hd__decap_4
X_0822_ PAR_IN2[17] _0956_/B _0822_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0801__A PAR_IN2[25] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_3 VSS VDD sky130_fd_sc_hd__decap_6
X_0684_ _0831_/A _0684_/B _0684_/C _0684_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0520__B _0519_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0753_ PAR_IN1[21] _0741_/B _0753_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0853__A2 _0637_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_297 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0711__A _0831_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_64 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_52 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_41 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_7_202 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_253 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_264 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_84 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0621__A _0618_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0532__A1 _0559_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_150 VSS VDD sky130_fd_sc_hd__decap_3
X_1021_ _1021_/D COUNT[2] RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_0805_ PAR_IN4[25] _0730_/X _0732_/X _0805_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0771__A1 PAR_IN7[29] VSS VDD sky130_fd_sc_hd__diode_2
X_0736_ PAR_IN7[11] _0706_/X _0735_/X _0736_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0531__A INTERNAL_FINISH VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0888__D _0887_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0598_ _0603_/A SAMPLE_COUNT[0] _0603_/C _0618_/B _0599_/A VSS VDD sky130_fd_sc_hd__and4_4
X_0667_ _0809_/A _0683_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_29_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_186 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_120 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0706__A _0705_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0826__A2 _0692_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1003__A2 _0597_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_54 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_21 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_10 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_52 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_164 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_153 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_109 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0616__A _0792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_194 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_384 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ COUNT[5] _0521_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_3_293 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_172 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_131 VSS VDD sky130_fd_sc_hd__fill_2
X_1004_ PAR_IN3[20] _0724_/A _1004_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0526__A _0603_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0899__C _0898_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0992__A1 PAR_IN8[4] VSS VDD sky130_fd_sc_hd__diode_2
X_0719_ PAR_IN8[27] _0657_/X _0718_/X _0719_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_25_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_167 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_87 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_75 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_123 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_170 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_131 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_186 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0974__A1 PAR_IN8[28] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_181 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_201 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_278 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_39_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_167 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0717__A1 PAR_IN4[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_292 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_259 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_105 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_13_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_138 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_149 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0708__A1 PAR_IN7[19] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_218 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_226 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_215 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0892__B1 _0891_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0984_ PAR_IN7[12] _0705_/X _0983_/X _0984_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_44_292 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0644__B1 _0643_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0947__A1 PAR_IN3[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_226 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_207 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0938__A1 PAR_IN8[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_126 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_148 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_44 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_74 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0874__B1 _0590_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0624__A PAR_IN7[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_292 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0929__A1 PAR_IN4[0] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0997__C _0996_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_130 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0617__B1 _0616_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0518__B _0517_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_270 VSS VDD sky130_fd_sc_hd__decap_4
X_0967_ PAR_IN1[28] _0967_/B _0967_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_32_284 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0534__A _0562_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0898_ _0898_/A _0898_/B _0898_/C _0897_/X _0898_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0709__A _0700_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1027__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0619__A _0619_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_47 VSS VDD sky130_fd_sc_hd__decap_12
X_0752_ _0512_/X _0741_/X _0751_/X _0752_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0821_ PAR_IN1[17] _0593_/B _0821_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0801__B _0956_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_3 VSS VDD sky130_fd_sc_hd__decap_3
X_0683_ _0683_/A _0668_/X _0683_/C _0684_/C VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_49_192 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0838__B1 _0837_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0529__A _0552_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0711__B _0711_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0902__A PAR_IN4[22] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_221 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_52 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_258 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0621__B _0581_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1020_ _1020_/D COUNT[1] RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0532__A2 _0531_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_173 VSS VDD sky130_fd_sc_hd__decap_6
X_0804_ PAR_IN8[25] _0676_/X _0803_/X _0804_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0812__A PAR_IN2[1] VSS VDD sky130_fd_sc_hd__diode_2
X_0735_ PAR_IN6[11] _0744_/B _0735_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0597_ _0994_/B _0597_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0771__A2 _0706_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0666_ _0627_/A _0666_/B _0665_/X _0684_/B VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_52_132 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_110 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_198 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0722__A _0593_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_140 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_352 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_52 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_30 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_330 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_162 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_385 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0632__A PAR_IN1[31] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_13 VSS VDD sky130_fd_sc_hd__fill_2
X_0520_ _0810_/A _0519_/X _0520_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_3_272 VSS VDD sky130_fd_sc_hd__fill_2
X_1003_ PAR_IN6[20] _0597_/X _0616_/X _1003_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_19_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_198 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0542__A SAMPLE_COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0992__A2 _0676_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0718_ PAR_IN5[27] _0694_/B _0718_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0649_ PAR_IN7[31] _0645_/X _0648_/X _0649_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_40_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_22 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_253 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_0_231 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_257 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_235 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0627__A _0627_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_146 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_160 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0974__A2 _0676_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_235 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0537__A SAMPLE_COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0717__A2 _0642_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_65 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_102 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0910__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0708__A2 _0706_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0892__A1 PAR_IN6[14] VSS VDD sky130_fd_sc_hd__diode_2
X_0983_ PAR_IN6[12] _0994_/B _0983_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0947__A2 _0634_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_172 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0644__A1 PAR_IN4[31] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_190 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0820__A _0627_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_282 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0730__A _0787_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0938__A2 _0657_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_12 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1023__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_86 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_238 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0874__A1 PAR_IN3[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_63 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0929__A2 _0600_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0624__B _0645_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0640__A PAR_IN5[31] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_142 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_175 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0617__A1 PAR_IN3[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_219 VSS VDD sky130_fd_sc_hd__fill_2
X_0966_ COUNT[2] _0944_/Y _0965_/Y _0966_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0897_ PAR_IN2[14] _0925_/B _0896_/X _0897_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0550__A _0577_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_90 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0709__B _0709_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0725__A _0724_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_263 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_23_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_23_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_189 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_167 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_15 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0635__A _0634_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_59 VSS VDD sky130_fd_sc_hd__decap_3
X_0820_ _0627_/A _0811_/X _0819_/X _0820_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0751_ _0751_/A _0745_/X _0751_/C _0750_/X _0751_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_9_46 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_285 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_3 VSS VDD sky130_fd_sc_hd__decap_3
X_0682_ _0682_/A _0674_/X _0675_/X _0682_/D _0683_/C VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_49_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_37_300 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0838__A1 PAR_IN2[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_266 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_255 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0545__A _0586_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0949_ PAR_IN7[24] _0705_/X _0948_/X _0953_/B VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0711__C _0711_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_32 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0902__B _0870_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_233 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0621__C _0603_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_8 VSS VDD sky130_fd_sc_hd__fill_2
X_0803_ PAR_IN5[25] _0803_/B _0803_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0812__B _0956_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0665_ _0665_/A _0659_/X _0660_/X _0664_/X _0665_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0734_ PAR_IN4[11] _0731_/X _0733_/X _0734_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_6_292 VSS VDD sky130_fd_sc_hd__decap_4
X_0596_ _0862_/B _0994_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_29_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_130 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0995__B1 _0994_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_78 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_207 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_152 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_386 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_111 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_320 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0913__A PAR_IN5[6] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0632__B _0631_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_25 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_6_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_122 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_152 VSS VDD sky130_fd_sc_hd__fill_1
X_1002_ PAR_IN2[20] _0620_/X _1001_/X _1002_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0729__B1 _0728_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0648_ PAR_IN6[31] _0673_/B _0648_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0717_ PAR_IN4[27] _0642_/X _0643_/X _0717_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0579_ _0559_/X _0524_/Y _0578_/X _1023_/D VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__0733__A _0732_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_199 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_111 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_12 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_225 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_0_265 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0627__B _0593_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0959__B1 _0958_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0643__A _0792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_103 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_150 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_199 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_158 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0553__A _0581_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_239 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_291 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_280 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0728__A PAR_IN5[11] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_261 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_87 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_54 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_99 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_114 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0910__B _0901_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0638__A PAR_IN2[31] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_272 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0644__A2 _0642_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0892__A2 _0646_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0982_ PAR_IN4[12] _0730_/X _0732_/X _0982_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_8_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_195 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0820__B _0811_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_297 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_231 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_294 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_106 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_139 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_7 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_21 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_206 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_231 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0874__A2 _0634_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_75 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0640__B _0610_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_154 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0617__A2 _0614_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_283 VSS VDD sky130_fd_sc_hd__fill_2
X_0965_ _0965_/A _0954_/X _0964_/X _0965_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0896_ PAR_IN7[14] _0896_/B _0896_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0831__A _0831_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_231 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0709__C _0703_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_209 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0741__A PAR_IN1[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_275 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_23_56 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_124 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_86 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_27 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0916__A PAR_IN7[6] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_58 VSS VDD sky130_fd_sc_hd__decap_3
X_0750_ PAR_IN8[5] _0677_/X _0749_/X _0750_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0681_ PAR_IN8[23] _0677_/X _0680_/X _0682_/D VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0651__A _0809_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_29_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_172 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0838__A2 _0637_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0948_ PAR_IN6[24] _0662_/A _0948_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0561__A _0573_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_212 VSS VDD sky130_fd_sc_hd__fill_2
X_0879_ _0944_/A _0879_/B _0879_/C _0879_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_47_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_23 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_34_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_32 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0621__D _0621_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_197 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_186 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_142 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_301 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0646__A _0595_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0802_ PAR_IN3[25] _0724_/X _0801_/X _0808_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0664_ PAR_IN7[7] _0645_/X _0663_/X _0664_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0733_ _0732_/X _0733_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0595_ _0595_/A _0862_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_40_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_37_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_164 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0995__A1 PAR_IN7[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_68 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_21 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_120 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_304 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_387 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_98 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_332 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_145 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_321 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0913__B _0747_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_7 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_3_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_90 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0674__B1 _0673_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_307 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_197 VSS VDD sky130_fd_sc_hd__fill_2
X_1001_ PAR_IN8[20] _0656_/A _1001_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0729__A1 PAR_IN8[11] VSS VDD sky130_fd_sc_hd__diode_2
X_0578_ _0512_/X _0577_/X _0562_/X _0578_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0647_ _0646_/X _0673_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0716_ PAR_IN7[27] _0645_/X _0715_/X _0720_/B VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_25_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_204 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_0_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_222 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0924__A PAR_IN1[0] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0627__C _0626_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0959__A1 PAR_IN8[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_137 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_140 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_3 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0895__B1 _0590_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_104 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0553__B _0581_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_91 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_273 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0744__A PAR_IN6[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_23 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0728__B _0694_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_148 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0910__C _0910_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_229 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_207 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_49 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0638__B _0699_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0981_ PAR_IN8[12] _0657_/A _0980_/X _0985_/B VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0654__A PAR_IN2[7] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0820__C _0819_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_181 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0829__A _0823_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_276 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_118 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_33 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0739__A _0965_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_229 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_87 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_284 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_41_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_310 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_199 VSS VDD sky130_fd_sc_hd__fill_2
X_0964_ _0627_/A _0955_/X _0963_/X _0964_/X VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_32_298 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_276 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_295 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0831__B _0820_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0895_ PAR_IN3[14] _0634_/A _0590_/A _0898_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0709__D _0708_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0559__A _0559_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_254 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0741__B _0741_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_76 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0916__B _0623_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0932__A _0932_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_15 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_298 VSS VDD sky130_fd_sc_hd__fill_1
X_0680_ PAR_IN5[23] _0694_/B _0680_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0651__B _0651_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_184 VSS VDD sky130_fd_sc_hd__fill_2
X_0947_ PAR_IN3[24] _0634_/X _0946_/X _0953_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0842__A PAR_IN3[10] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0561__B _0560_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_280 VSS VDD sky130_fd_sc_hd__fill_1
X_0878_ _0510_/X _0869_/X _0878_/C _0879_/C VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0752__A _0512_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_257 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_165 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_305 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0927__A PAR_IN6[0] VSS VDD sky130_fd_sc_hd__diode_2
X_0801_ PAR_IN2[25] _0956_/B _0801_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0662__A _0662_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0663_ PAR_IN6[7] _0744_/B _0663_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_41_3 VSS VDD sky130_fd_sc_hd__decap_3
X_0732_ _0792_/A _0732_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_6_261 VSS VDD sky130_fd_sc_hd__fill_2
X_0594_ _0603_/C SAMPLE_COUNT[2] _0618_/C _0603_/B _0595_/A VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__0837__A PAR_IN4[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_82 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_135 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_102 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0995__A2 _0689_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_14 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_12 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_102 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_300 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0747__A _0747_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_316 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_377 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1020__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0657__A _0657_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_110 VSS VDD sky130_fd_sc_hd__fill_1
X_1000_ PAR_IN5[20] _0749_/B _0999_/X _1000_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_13_7 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0674__A1 PAR_IN7[23] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_135 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_113 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0729__A2 _0657_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0715_ PAR_IN6[27] _0673_/B _0715_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0577_ _0577_/A _0520_/X _0577_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0646_ _0595_/A _0646_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_25_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_57 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1026__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_249 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0924__B _0924_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_130 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__A2 _0676_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0940__A PAR_IN6[16] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_163 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_205 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0895__A1 PAR_IN3[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_182 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1011__A COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_138 VSS VDD sky130_fd_sc_hd__decap_12
X_0629_ _0976_/A _0809_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_53_230 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0744__B _0744_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_260 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_46 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_171 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0935__A PAR_IN2[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_271 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_252 VSS VDD sky130_fd_sc_hd__decap_12
X_0980_ PAR_IN5[12] _0930_/B _0980_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0654__B _0699_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_160 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0670__A _0946_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1006__A _1000_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0829__B _0829_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0845__A _0510_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_244 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0580__A _0550_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_307 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0556__B1 _0533_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_89 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0739__B _0739_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_44 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_299 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_41_200 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_241 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0795__B1 _0794_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_134 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0665__A _0665_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_252 VSS VDD sky130_fd_sc_hd__fill_2
X_0963_ _0957_/X _0959_/X _0963_/C _0962_/X _0963_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0831__C _0831_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0894_ PAR_IN8[14] _0907_/B _0893_/X _0898_/B VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_4_93 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_11 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0932__B _0928_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0651__C _0650_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0768__B1 _0767_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_288 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_196 VSS VDD sky130_fd_sc_hd__fill_1
X_0946_ PAR_IN2[24] _0946_/B _0946_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0842__B _0842_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_247 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_225 VSS VDD sky130_fd_sc_hd__fill_2
X_0877_ _0871_/X _0873_/X _0877_/C _0876_/X _0878_/C VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0931__B1 _0930_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_23 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0752__B _0741_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_3 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0922__B1 _0900_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0927__B _0646_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0943__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_317 VSS VDD sky130_fd_sc_hd__fill_2
X_0731_ _0730_/X _0731_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_24_90 VSS VDD sky130_fd_sc_hd__fill_2
X_0800_ _0619_/A _0956_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0593_ PAR_IN1[15] _0593_/B _0593_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0662_ _0662_/A _0744_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_34_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_284 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0837__B _0599_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_100 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_158 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_147 VSS VDD sky130_fd_sc_hd__decap_6
X_0929_ PAR_IN4[0] _0600_/X _0792_/X _0929_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_45_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_34 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_334 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__A _0831_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_378 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_254 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_133 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0673__A PAR_IN6[23] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0674__A2 _0645_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_158 VSS VDD sky130_fd_sc_hd__fill_2
X_0645_ _0645_/A _0645_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0714_ PAR_IN3[27] _0635_/X _0713_/X _0714_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1009__A _1009_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0576_ _0559_/X _0573_/Y _0575_/X _1022_/D VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__0583__A _0534_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_128 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_228 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_131 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_158 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0940__B _0662_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_186 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_239 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_217 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0668__A PAR_IN1[23] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0895__A2 _0634_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_250 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_0 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1011__B _0923_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0628_ COUNT[4] _0976_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_38_272 VSS VDD sky130_fd_sc_hd__decap_3
X_0559_ _0559_/A _0559_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_53_242 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_106 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_264 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0935__B _0946_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_250 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0951__A PAR_IN5[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_172 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_176 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1006__B _1002_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0829__C _0826_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_256 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0845__B _0836_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1016__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0580__B _0530_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0739__C _0738_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0556__A1 _0550_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_264 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_56 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_41_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_234 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0795__A1 PAR_IN2[9] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_146 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_157 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_179 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0946__A PAR_IN2[24] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0665__B _0659_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0962_ PAR_IN7[8] _0689_/X _0961_/X _0962_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0893_ PAR_IN5[14] _0608_/A _0893_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0856__A _0514_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0591__A _0591_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_278 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_48 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_256 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0932__C _0929_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0768__A1 PAR_IN8[29] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_8 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_307 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_49_142 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_171 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0676__A _0656_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_215 VSS VDD sky130_fd_sc_hd__decap_3
X_0945_ PAR_IN1[24] _0967_/B _0945_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0876_ PAR_IN2[2] _0637_/A _0875_/X _0876_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0931__A1 PAR_IN8[0] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0586__A _0586_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0695__B1 _0694_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0752__C _0751_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0922__A1 _0515_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0922__B2 _0921_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0943__B _0934_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0730_ _0787_/B _0730_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0661_ _0862_/B _0662_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_24_80 VSS VDD sky130_fd_sc_hd__decap_8
X_0592_ _0924_/B _0593_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_27_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_51 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_73 VSS VDD sky130_fd_sc_hd__fill_2
X_0928_ PAR_IN7[0] _0645_/A _0927_/X _0928_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0859_ _0599_/A _0870_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_45_13 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_36 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_181 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_368 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_68 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_335 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_115 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_324 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_178 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0763__B _0752_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_379 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0840__B1 _0839_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_222 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0954__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0659__B1 _0658_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_148 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_126 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_123 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0673__B _0673_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_90 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1009__B _0987_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0644_ PAR_IN4[31] _0642_/X _0643_/X _0644_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0713_ PAR_IN2[27] _0671_/B _0713_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0575_ _0577_/A _0965_/A _0562_/X _0575_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_33_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_159 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_115 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0583__B _0583_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_38 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_207 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_269 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0774__A PAR_IN1[13] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_104 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0813__B1 _0812_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_107 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_132 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0668__B _0631_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0684__A _0831_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_1 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0804__B1 _0803_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_140 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1011__C _1010_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_181 VSS VDD sky130_fd_sc_hd__fill_2
X_0627_ _0627_/A _0593_/X _0626_/X _0627_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0558_ _0559_/A COUNT[0] _0557_/X _0535_/X _0534_/X _0558_/Y VSS VDD sky130_fd_sc_hd__a2111oi_4
XANTENNA__0859__A _0599_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_15 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0594__A _0603_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_36 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_14 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_276 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_262 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0951__B _0803_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_144 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_12_140 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_184 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0679__A _0930_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_199 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_221 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1006__C _1003_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0829__D _0829_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_268 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_202 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0845__C _0844_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0580__C COUNT[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0556__A2 _0554_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0589__A _0615_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_47 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0795__A2 _0620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_114 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0946__B _0946_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_221 VSS VDD sky130_fd_sc_hd__fill_2
X_0961_ PAR_IN6[8] _0994_/B _0961_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0665__C _0660_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_257 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_32_235 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_243 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_290 VSS VDD sky130_fd_sc_hd__decap_12
X_0892_ PAR_IN6[14] _0646_/X _0891_/X _0898_/A VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_4_180 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0856__B _0845_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0872__A PAR_IN5[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_316 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0782__A _0782_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_235 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_246 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0932__D _0931_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0768__A2 _0677_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_176 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0692__A _0787_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0944_ _0944_/A _0933_/X _0943_/X _0944_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0875_ PAR_IN7[2] _0896_/B _0875_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_9_283 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0931__A2 _0657_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0695__A1 PAR_IN8[3] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0867__A _0867_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0586__B _0586_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_69 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_11_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0777__A PAR_IN6[13] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0922__A2 _0856_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_179 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0943__C _0942_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0591_ _0591_/A _0924_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0660_ PAR_IN4[7] _0642_/X _0643_/X _0660_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_10_282 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_293 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_30 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0687__A PAR_IN2[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_190 VSS VDD sky130_fd_sc_hd__decap_4
X_0927_ PAR_IN6[0] _0646_/X _0927_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0597__A _0994_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0858_ PAR_IN1[18] _0901_/B _0868_/B VSS VDD sky130_fd_sc_hd__or2_4
X_0789_ _0608_/A _0789_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_28_135 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_369 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_127 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_325 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0840__A1 PAR_IN7[10] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0763__C _0763_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_102 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_3_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_61 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0954__B _0945_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0659__A1 PAR_IN8[7] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0970__A PAR_IN6[28] VSS VDD sky130_fd_sc_hd__diode_2
X_0574_ _0810_/A _0965_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1009__C _1009_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0643_ _0792_/A _0643_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0712_ PAR_IN1[27] _0631_/X _0721_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_25_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0880__A PAR_IN1[30] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_215 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_100 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0774__B _0741_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0813__A1 PAR_IN3[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_193 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_182 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_199 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0790__A PAR_IN5[9] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_144 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_71 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_263 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0965__A _0965_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0804__A1 PAR_IN8[25] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_296 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0684__B _0684_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_119 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_2 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_160 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0568__B1 _0562_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_62 VSS VDD sky130_fd_sc_hd__fill_2
X_0626_ _0626_/A _0611_/X _0617_/X _0625_/X _0626_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0557_ _0577_/A COUNT[5] _0518_/A _0557_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_53_211 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0875__A PAR_IN7[2] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0594__B SAMPLE_COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_29_241 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0785__A _1009_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_233 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1006__D _1006_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_247 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0580__D _0533_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_29 VSS VDD sky130_fd_sc_hd__fill_2
X_0609_ _0747_/A _0610_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_41_225 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_41_203 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_303 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0952__B1 _0951_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_310 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0665__D _0664_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_81 VSS VDD sky130_fd_sc_hd__fill_2
X_0960_ PAR_IN4[8] _0692_/X _0732_/X _0963_/C VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_32_269 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_299 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_266 VSS VDD sky130_fd_sc_hd__fill_2
X_0891_ PAR_IN4[14] _0870_/B _0891_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0856__C _0855_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_203 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0872__B _0608_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_39 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_28 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0782__B _0778_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_83 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_155 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1023__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_195 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_91 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0973__A PAR_IN5[28] VSS VDD sky130_fd_sc_hd__diode_2
X_0943_ _0976_/A _0934_/X _0942_/X _0943_/X VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_9_240 VSS VDD sky130_fd_sc_hd__decap_4
X_0874_ PAR_IN3[2] _0634_/A _0590_/A _0877_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0695__A2 _0657_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0867__B _0863_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0586__C _0618_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_38 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0883__A PAR_IN6[30] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0777__B _0597_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0922__A3 _0879_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_103 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_24_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_60 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0968__A PAR_IN2[28] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_70 VSS VDD sky130_fd_sc_hd__decap_4
X_0590_ _0590_/A _0591_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_6_276 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_6_265 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0687__B _0699_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_106 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_86 VSS VDD sky130_fd_sc_hd__decap_12
X_0926_ PAR_IN3[0] _0634_/X _0925_/X _0932_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0857_ _0591_/A _0901_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_20_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_18 VSS VDD sky130_fd_sc_hd__fill_1
X_0788_ PAR_IN6[9] _0744_/B _0787_/X _0788_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0878__A _0510_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_48 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_26 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_158 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_359 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_191 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0840__A2 _0623_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_268 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_213 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_73 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0659__A2 _0657_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0954__C _0953_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_80 VSS VDD sky130_fd_sc_hd__fill_2
X_0711_ _0831_/A _0711_/B _0711_/C _0740_/B VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0970__B _0646_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0642_ _0600_/X _0642_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_32_3 VSS VDD sky130_fd_sc_hd__fill_2
X_0573_ _0573_/A _0573_/B _0573_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__0698__A PAR_IN1[19] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_106 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1019__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_172 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_18 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0880__B _0901_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0909_ _0909_/A _0905_/X _0909_/C _0908_/X _0910_/C VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_0_249 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_101 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_134 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0813__A2 _0614_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0790__B _0789_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_145 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_220 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0965__B _0954_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0684__C _0684_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0804__A2 _0676_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_91 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_3 VSS VDD sky130_fd_sc_hd__decap_3
X_0625_ PAR_IN2[15] _0620_/X _0624_/X _0625_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_30_186 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0568__A1 _0550_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0556_ _0550_/X _0554_/X _0533_/A _0556_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_38_297 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0875__B _0896_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0594__C _0618_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0891__A PAR_IN4[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_164 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_142 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_275 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0785__B _0763_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_245 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_164 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0976__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_278 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1022__D _1022_/D VSS VDD sky130_fd_sc_hd__diode_2
X_0608_ _0608_/A _0747_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0886__A PAR_IN8[30] VSS VDD sky130_fd_sc_hd__diode_2
X_0539_ _0535_/X _0536_/X _0621_/D _0540_/C VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_53_15 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_256 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_138 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0796__A _0788_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0952__A1 PAR_IN8[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_81 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_270 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_215 VSS VDD sky130_fd_sc_hd__fill_2
X_0890_ PAR_IN1[14] _0901_/B _0899_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_4_42 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1017__D _1017_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_215 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_270 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0782__C _0779_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0973__B _0803_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0861__B1 _0860_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0942_ _0936_/X _0938_/X _0939_/X _0941_/X _0942_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_20_229 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_207 VSS VDD sky130_fd_sc_hd__decap_3
X_0873_ PAR_IN8[2] _0907_/B _0872_/X _0873_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_13_281 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0867__C _0864_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_307 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0883__B _0862_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_159 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_137 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0843__B1 _0842_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_233 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_40_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0968__B _0925_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_7 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_148 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_104 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_98 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_170 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0834__B1 _0785_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0787_ PAR_IN4[9] _0787_/B _0787_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0925_ PAR_IN2[0] _0925_/B _0925_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0856_ _0514_/A _0845_/X _0855_/X _0856_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_29_17 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0878__B _0869_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_316 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_170 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_310 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0825__B1 _0824_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_151 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_349 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_236 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1002__B1 _1001_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_85 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_148 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_94 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_173 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0816__B1 _0616_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_107 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_310 VSS VDD sky130_fd_sc_hd__decap_8
X_0710_ _0683_/A _0710_/B _0709_/X _0711_/C VSS VDD sky130_fd_sc_hd__and3_4
X_0641_ PAR_IN8[31] _0606_/X _0640_/X _0650_/B VSS VDD sky130_fd_sc_hd__a21o_4
X_0572_ _0831_/A _0566_/Y _0520_/X _0573_/B VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_25_3 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0698__B _0631_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1025__D _0540_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0807__B1 _0806_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_151 VSS VDD sky130_fd_sc_hd__decap_4
X_0908_ PAR_IN2[22] _0956_/B _0907_/X _0908_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0889__A COUNT[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_228 VSS VDD sky130_fd_sc_hd__fill_1
X_0839_ PAR_IN6[10] _0595_/A _0839_/X VSS VDD sky130_fd_sc_hd__and2_4
XPHY_102 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_135 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0799__A PAR_IN1[25] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_317 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_168 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_232 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_81 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0965__C _0964_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_154 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_4 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_184 VSS VDD sky130_fd_sc_hd__fill_2
X_0624_ PAR_IN7[15] _0645_/A _0624_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0568__A2 _1009_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_243 VSS VDD sky130_fd_sc_hd__fill_2
X_0555_ _0550_/X _0530_/D _0534_/X _0553_/Y _0554_/X _0555_/Y VSS VDD sky130_fd_sc_hd__a2111oi_4
XFILLER_38_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_276 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0594__D _0603_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0891__B _0870_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_287 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_29_254 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0785__C _0785_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_268 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1017__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_40 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_147 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_198 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0976__B _0967_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_213 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_202 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0886__B _0852_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0538_ _0586_/B _0621_/D VSS VDD sky130_fd_sc_hd__buf_1
X_0607_ _0618_/A _0581_/B _0618_/C _0621_/D _0608_/A VSS VDD sky130_fd_sc_hd__and4_4
XFILLER_37_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_268 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0796__B _0791_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0952__A2 _0606_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_205 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_72 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_71 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_260 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_249 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_25_290 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0987__A _0810_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_172 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_290 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_109 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_308 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0782__D _0782_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_293 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_30 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0600__A _0787_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_131 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_49_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_164 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_175 VSS VDD sky130_fd_sc_hd__decap_8
X_0941_ PAR_IN7[16] _0705_/X _0940_/X _0941_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0861__A1 PAR_IN5[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_253 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_9_297 VSS VDD sky130_fd_sc_hd__fill_2
X_0872_ PAR_IN5[2] _0608_/A _0872_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_13_293 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0510__A _0509_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0867__D _0866_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1028__D _0556_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_311 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0843__A1 PAR_IN5[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_40 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_70 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_92 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_66 VSS VDD sky130_fd_sc_hd__fill_1
X_0924_ PAR_IN1[0] _0924_/B _0924_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_45_182 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0834__B2 _0833_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0834__A1 _0517_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0786_ PAR_IN1[9] _0967_/B _0786_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0855_ COUNT[4] _0846_/X _0854_/X _0855_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0878__C _0878_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_116 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0522__B1 _0521_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_339 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_119 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_328 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0825__A1 PAR_IN8[17] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1002__A1 PAR_IN2[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0816__A1 PAR_IN4[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_94 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_50 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_182 VSS VDD sky130_fd_sc_hd__fill_1
X_0571_ _0944_/A _0831_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0640_ PAR_IN5[31] _0610_/B _0640_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_18_3 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0807__A1 PAR_IN7[25] VSS VDD sky130_fd_sc_hd__diode_2
X_0907_ PAR_IN8[22] _0907_/B _0907_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0838_ PAR_IN2[10] _0637_/A _0837_/X _0838_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0743__B1 _0742_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_218 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_207 VSS VDD sky130_fd_sc_hd__decap_8
X_0769_ PAR_IN4[29] _0731_/X _0733_/X _0772_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0889__B _0889_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_119 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_103 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_125 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0799__B _0988_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0982__B1 _0732_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_96 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_85 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0734__B1 _0733_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_93 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_5 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_130 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_174 VSS VDD sky130_fd_sc_hd__decap_4
X_0623_ _0623_/A _0645_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_87 VSS VDD sky130_fd_sc_hd__fill_2
X_0554_ _0581_/B _0581_/D _0554_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_38_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_42_18 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_100 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_200 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0716__B1 _0715_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_280 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_8_104 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_177 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0603__A _0603_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0976__C _0976_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_236 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_225 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0513__A COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_192 VSS VDD sky130_fd_sc_hd__fill_2
X_0537_ SAMPLE_COUNT[0] _0586_/B VSS VDD sky130_fd_sc_hd__inv_8
X_0606_ _0656_/A _0606_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_37_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_203 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_291 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_118 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0796__C _0796_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_203 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_225 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0928__B1 _0927_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0987__B _0976_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_140 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_66 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0508__A SAMPLE_COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_250 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0919__B1 _0509_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_53 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_83 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_61 VSS VDD sky130_fd_sc_hd__decap_4
X_0940_ PAR_IN6[16] _0662_/A _0940_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0861__A2 _0789_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_221 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0998__A PAR_IN1[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_276 VSS VDD sky130_fd_sc_hd__decap_4
X_0871_ PAR_IN6[2] _0646_/X _0870_/X _0871_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_48_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_19 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_209 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0701__A PAR_IN5[19] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0843__A2 _0789_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_257 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_194 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_117 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_301 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0834__A2 _0685_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_34 VSS VDD sky130_fd_sc_hd__fill_2
X_0854_ _0848_/X _0854_/B _0851_/X _0853_/X _0854_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0923_ COUNT[1] _0922_/X _0923_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0785_ _1009_/A _0763_/Y _0785_/C _0785_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0521__A COUNT[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_290 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0522__A1 _0512_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_131 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_329 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0825__A2 _0606_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1002__A2 _0620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_43 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0816__A2 _0692_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_172 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_117 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_74 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_142 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_62 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0606__A _0656_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_94 VSS VDD sky130_fd_sc_hd__decap_4
X_0570_ COUNT[3] _0944_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0807__A2 _0689_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0516__A COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_194 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_150 VSS VDD sky130_fd_sc_hd__decap_3
X_0837_ PAR_IN4[10] _0599_/A _0837_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0906_ PAR_IN3[22] _0724_/A _0590_/A _0909_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0889__C _0889_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0699_ PAR_IN2[19] _0699_/B _0699_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0743__A1 PAR_IN3[5] VSS VDD sky130_fd_sc_hd__diode_2
X_0768_ PAR_IN8[29] _0677_/X _0767_/X _0768_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_24_120 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_104 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_175 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_126 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0982__A1 PAR_IN4[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_75 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_31 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0734__A1 PAR_IN4[11] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_267 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_6 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_3 VSS VDD sky130_fd_sc_hd__fill_2
X_0622_ _0896_/B _0623_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0553_ _0581_/B _0581_/D _0553_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_38_256 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0716__A1 PAR_IN7[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_248 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_75 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_74 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_32_41 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_116 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_138 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_112 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0603__B _0603_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1026__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_270 VSS VDD sky130_fd_sc_hd__decap_4
X_0605_ _0907_/B _0656_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0536_ _0559_/A _0573_/A _0536_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_26_215 VSS VDD sky130_fd_sc_hd__fill_2
X_1019_ _0558_/Y COUNT[0] RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0882__B1 _0881_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0704__A _0896_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0796__D _0795_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_237 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0625__B1 _0624_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_229 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_85 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0873__B1 _0872_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0928__A1 PAR_IN7[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_95 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0614__A _0724_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0987__C _0986_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_78 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_23_218 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0864__B1 _0615_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_240 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0524__A _0573_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0919__A1 PAR_IN1[6] VSS VDD sky130_fd_sc_hd__diode_2
X_0519_ _0515_/Y _0519_/B _0519_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_13_10 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_87 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_104 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_144 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_159 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_310 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0609__A _0747_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0870_ PAR_IN4[2] _0870_/B _0870_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_9_200 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_240 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0998__B _0593_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0519__A _0515_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_19 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1014__B1 _1013_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0999_ PAR_IN7[20] _0794_/B _0999_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0701__B _0694_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_107 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_310 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0828__B1 _0827_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_74 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_63 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_41 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1005__B1 _1004_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_247 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_276 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_184 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0834__A3 _0740_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0853_ PAR_IN2[26] _0637_/A _0852_/X _0853_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0922_ _0515_/Y _0856_/X _0879_/X _0900_/X _0921_/X _0922_/X VSS VDD sky130_fd_sc_hd__a32o_4
X_0784_ _0965_/A _0784_/B _0783_/X _0785_/C VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_28_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0522__A2 _0520_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_198 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_165 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_319 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0712__A PAR_IN1[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_129 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_74 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_184 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_86 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_165 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_305 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0622__A _0896_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_272 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_110 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_184 VSS VDD sky130_fd_sc_hd__decap_4
X_0836_ PAR_IN1[10] _0591_/A _0836_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0905_ PAR_IN7[22] _0794_/B _0904_/X _0905_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0767_ PAR_IN5[29] _0749_/B _0767_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0743__A2 _0725_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0698_ PAR_IN1[19] _0631_/X _0710_/B VSS VDD sky130_fd_sc_hd__or2_4
XPHY_105 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0707__A PAR_IN6[19] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_143 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_132 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_116 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_127 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_309 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_316 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0982__A2 _0730_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0734__A2 _0731_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_102 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_7 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_34 VSS VDD sky130_fd_sc_hd__fill_2
X_0621_ _0618_/A _0581_/B _0603_/A _0621_/D _0896_/B VSS VDD sky130_fd_sc_hd__and4_4
XFILLER_23_3 VSS VDD sky130_fd_sc_hd__fill_2
X_0552_ _0552_/A _0547_/B _0581_/D VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_53_249 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_268 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0527__A _0618_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_168 VSS VDD sky130_fd_sc_hd__fill_1
X_0819_ _0819_/A _0815_/X _0816_/X _0818_/X _0819_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0716__A2 _0645_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_279 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_86 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0603__C _0603_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0900__A _0810_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_219 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_208 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0810__A _0810_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0604_ _0852_/B _0907_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_161 VSS VDD sky130_fd_sc_hd__decap_4
X_0535_ COMPLETE _0535_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0882__A1 PAR_IN5[30] VSS VDD sky130_fd_sc_hd__diode_2
X_1018_ _0581_/X COMPLETE RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0720__A _0714_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_53 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_249 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0873__A1 PAR_IN8[2] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0625__A1 PAR_IN2[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_85 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_219 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_97 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0928__A2 _0645_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0630__A _0924_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1022__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0864__A1 PAR_IN3[18] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0919__A2 _0924_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0518_ _0518_/A _0517_/Y _0519_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0540__A _0530_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_285 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_263 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0715__A PAR_IN6[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_219 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_77 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0791__B1 _0790_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_138 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_123 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_263 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_285 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_300 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0519__B _0519_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0535__A COMPLETE VSS VDD sky130_fd_sc_hd__diode_2
X_0998_ PAR_IN1[20] _0593_/B _1007_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1014__A1 _0535_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_119 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0828__A1 PAR_IN7[17] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_255 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1005__A1 PAR_IN4[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_174 VSS VDD sky130_fd_sc_hd__fill_2
X_0921_ _0910_/X _0920_/X COUNT[2] _0921_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_53_3 VSS VDD sky130_fd_sc_hd__decap_12
X_0852_ PAR_IN8[26] _0852_/B _0852_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0783_ _0512_/X _0783_/B _0783_/C _0783_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0755__B1 _0754_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_100 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_174 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_163 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_177 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_309 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0746__B1 _0733_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_218 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0712__B _0631_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_43 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_10 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_177 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_86 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_196 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_174 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_188 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_306 VSS VDD sky130_fd_sc_hd__decap_12
X_0904_ PAR_IN6[22] _0862_/B _0904_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0835_ COUNT[0] _0834_/Y _0835_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0697_ _0627_/A _0697_/B _0697_/C _0711_/B VSS VDD sky130_fd_sc_hd__and3_4
X_0766_ PAR_IN3[29] _0725_/X _0765_/X _0766_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0707__B _0744_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_106 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_128 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0723__A PAR_IN1[11] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0719__B1 _0718_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_258 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_85 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_46_41 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_169 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0633__A _0842_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_8 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_188 VSS VDD sky130_fd_sc_hd__decap_12
X_0620_ _0925_/B _0620_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_310 VSS VDD sky130_fd_sc_hd__decap_8
X_0551_ SAMPLE_COUNT[2] _0581_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_38_203 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0808__A _0808_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_291 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_247 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0949__B1 _0948_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_114 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0543__A _0603_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0818_ PAR_IN8[1] _0606_/X _0817_/X _0818_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0749_ PAR_IN5[5] _0749_/B _0749_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_44_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0718__A PAR_IN5[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_21 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_125 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_32 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_180 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0603__D SAMPLE_COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0900__B _0900_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0628__A COUNT[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_280 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_140 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0810__B _0810_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0534_ _0562_/B _0534_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_184 VSS VDD sky130_fd_sc_hd__fill_2
X_0603_ _0603_/A _0603_/B _0603_/C SAMPLE_COUNT[2] _0852_/B VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__0538__A _0586_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_261 VSS VDD sky130_fd_sc_hd__decap_12
X_1017_ _1017_/D INTERNAL_FINISH RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0882__A2 _0789_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0720__B _0720_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0555__D1 _0554_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_209 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_217 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0873__A2 _0907_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0625__A2 _0620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_42 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_294 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0911__A PAR_IN4[6] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_176 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_36 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0864__A2 _0634_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_261 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_275 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0821__A PAR_IN1[17] VSS VDD sky130_fd_sc_hd__diode_2
X_0517_ COUNT[1] _0517_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__0540__B _0534_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0715__B _0673_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_34 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0791__A1 PAR_IN8[9] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0731__A _0730_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_102 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_168 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_312 VSS VDD sky130_fd_sc_hd__decap_6
X_0997_ _0933_/A _0988_/X _0996_/X _0997_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1014__A2 SERIAL_OUT VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0551__A SAMPLE_COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_161 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_150 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_172 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0828__A2 _0689_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0726__A PAR_IN2[11] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1005__A2 _0692_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_74 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_153 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_15 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_197 VSS VDD sky130_fd_sc_hd__fill_2
X_0920_ _0918_/X _0919_/X _0944_/A _0920_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0636__A _0619_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0851_ PAR_IN3[26] _0842_/B _0615_/A _0851_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0782_ _0782_/A _0778_/X _0779_/X _0782_/D _0783_/C VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0755__A1 PAR_IN3[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_3 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_145 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0691__B1 _0690_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0746__A1 PAR_IN4[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_131 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_54 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_43 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_164 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_285 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_241 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_123 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_142 VSS VDD sky130_fd_sc_hd__decap_8
X_0903_ PAR_IN5[22] _0789_/X _0902_/X _0909_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0834_ _0517_/Y _0685_/Y _0740_/Y _0785_/Y _0833_/X _0834_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XFILLER_21_318 VSS VDD sky130_fd_sc_hd__fill_1
X_0765_ PAR_IN2[29] _0620_/X _0765_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0696_ _0688_/X _0691_/X _0696_/C _0695_/X _0697_/C VSS VDD sky130_fd_sc_hd__or4_4
XPHY_107 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0664__B1 _0663_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_178 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_129 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0723__B _0741_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_67 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0719__A1 PAR_IN8[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_64 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0655__B1 _0654_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_9 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_134 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_148 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_126 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_178 VSS VDD sky130_fd_sc_hd__fill_1
X_0550_ _0577_/A _0550_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_215 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0894__B1 _0893_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_218 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_53_207 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0808__B _0804_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_281 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0824__A PAR_IN5[17] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0949__A1 PAR_IN7[24] VSS VDD sky130_fd_sc_hd__diode_2
X_0817_ PAR_IN5[1] _0610_/B _0817_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0543__B _0603_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0679_ _0930_/B _0694_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0748_ _0803_/B _0749_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_29_237 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_204 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0718__B _0694_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0885__B1 _0590_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_295 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_32_11 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0900__C _0900_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0909__A _0909_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0876__B1 _0875_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_262 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_170 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0810__C _0809_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0602_ PAR_IN6[15] _0597_/X _0601_/X _0626_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0533_ _0533_/A _0562_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_7_196 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0819__A _0819_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_229 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_251 VSS VDD sky130_fd_sc_hd__decap_4
X_1016_ _1015_/X SERIAL_OUT RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0554__A _0581_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0720__C _0717_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_11 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0555__C1 _0553_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_66 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_273 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_229 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_43_54 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_243 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0911__B _0787_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_15 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_210 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_273 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_290 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0821__B _0593_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0540__C _0540_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0516_ COUNT[0] _0518_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_22_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0791__A2 _0657_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_147 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_87 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_65 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_38_32 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_232 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_191 VSS VDD sky130_fd_sc_hd__fill_2
X_0996_ _0990_/X _0992_/X _0996_/C _0995_/X _0996_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0832__A COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_56 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0726__B _0671_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_66 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0742__A PAR_IN2[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_206 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_235 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_31 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0652__A _0965_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0850_ PAR_IN7[26] _0623_/A _0849_/X _0854_/B VSS VDD sky130_fd_sc_hd__a21o_4
X_0781_ PAR_IN8[13] _0677_/X _0780_/X _0782_/D VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0755__A2 _0725_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_36_110 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0827__A PAR_IN6[17] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0691__A1 PAR_IN7[3] VSS VDD sky130_fd_sc_hd__diode_2
X_0979_ PAR_IN3[12] _0724_/X _0978_/X _0985_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0562__A COMPLETE VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0746__A2 _0731_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_47 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_176 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0737__A _0737_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_146 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_135 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_297 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_264 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_157 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_165 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0647__A _0646_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0833_ COUNT[1] _0832_/Y _0833_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0902_ PAR_IN4[22] _0870_/B _0902_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0695_ PAR_IN8[3] _0657_/X _0694_/X _0695_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0764_ PAR_IN1[29] _0741_/B _0773_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0664__A1 PAR_IN7[7] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_124 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_108 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_308 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_35 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0719__A2 _0657_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_205 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0655__A1 PAR_IN3[7] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_102 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0930__A PAR_IN5[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1025__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0808__C _0805_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_260 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_227 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0894__A1 PAR_IN8[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_149 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_138 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0824__B _0610_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0949__A2 _0705_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0816_ PAR_IN4[1] _0692_/X _0616_/X _0816_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0747_ _0747_/A _0803_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1001__A PAR_IN8[20] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0543__C _0524_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_216 VSS VDD sky130_fd_sc_hd__fill_2
X_0678_ _0747_/A _0930_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0582__B1 _0530_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_241 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_282 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0885__A1 PAR_IN3[30] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_171 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_79 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0909__B _0905_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0876__A1 PAR_IN2[2] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0925__A PAR_IN2[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_285 VSS VDD sky130_fd_sc_hd__decap_4
X_0601_ PAR_IN4[15] _0600_/X _0601_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_7_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_175 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_193 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0819__B _0815_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0564__B1 _0563_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_3 VSS VDD sky130_fd_sc_hd__decap_3
X_0532_ _0559_/A _0531_/Y READY _0533_/A VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__0835__A COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
X_1015_ _0533_/A _1014_/X _1015_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0554__B _0581_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0570__A COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_91 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0720__D _0719_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0555__B1 _0534_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_34 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_23 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_99 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_266 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_101 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_134 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0546__B1 _0618_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_230 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_291 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_285 VSS VDD sky130_fd_sc_hd__decap_3
X_0515_ COUNT[2] _0515_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__0565__A _0515_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0776__B1 _0775_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_7 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_314 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0700__B1 _0699_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_204 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_211 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_255 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_306 VSS VDD sky130_fd_sc_hd__decap_12
X_0995_ PAR_IN7[4] _0689_/X _0994_/X _0995_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0832__B _0810_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0758__B1 _0733_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_70 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_24_24 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0742__B _0671_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_12 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_21 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0921__B1 COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0933__A _0933_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0652__B _0627_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0780_ PAR_IN5[13] _0749_/B _0780_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_14_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_262 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0912__B1 _0911_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0827__B _0673_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_169 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_114 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0979__B1 _0978_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_199 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1004__A PAR_IN3[20] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0691__A2 _0689_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0978_ PAR_IN2[12] _0946_/B _0978_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0562__B _0562_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0903__B1 _0902_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_12 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_111 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0737__B _0729_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_169 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0753__A PAR_IN1[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_232 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_9 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0663__A PAR_IN6[7] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_136 VSS VDD sky130_fd_sc_hd__fill_2
X_0901_ PAR_IN1[22] _0901_/B _0901_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0832_ COUNT[2] _0810_/Y _0831_/Y _0832_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0763_ _0831_/A _0752_/X _0763_/C _0763_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0694_ PAR_IN5[3] _0694_/B _0694_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_51_3 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0664__A2 _0645_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0573__A _0573_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_169 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_147 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_109 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_217 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0748__A _0803_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_77 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0655__A2 _0635_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0930__B _0930_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0808__D _0807_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0658__A PAR_IN5[7] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_239 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0894__A2 _0907_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1001__B _0656_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_180 VSS VDD sky130_fd_sc_hd__fill_2
X_0815_ PAR_IN7[1] _0705_/X _0814_/X _0815_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0746_ PAR_IN4[5] _0731_/X _0733_/X _0751_/C VSS VDD sky130_fd_sc_hd__a21o_4
X_0677_ _0676_/X _0677_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0885__A2 _0634_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0582__B2 _0531_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0582__A1 _0535_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_36 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_58 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0558__D1 _0534_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0909__C _0909_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0876__A2 _0637_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0925__B _0925_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_242 VSS VDD sky130_fd_sc_hd__fill_2
X_0600_ _0787_/B _0600_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_22_90 VSS VDD sky130_fd_sc_hd__fill_2
X_0531_ INTERNAL_FINISH _0531_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_7_165 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0819__C _0816_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0564__A1 _0559_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0835__B _0834_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1014_ _0535_/X SERIAL_OUT _1013_/Y _1014_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_34_297 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1012__A SAMPLE_COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
X_0729_ PAR_IN8[11] _0657_/X _0728_/X _0729_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0555__A1 _0550_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_223 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_264 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0761__A _0761_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_168 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0546__A1 _0621_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_242 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_253 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_292 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_270 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0671__A PAR_IN2[23] VSS VDD sky130_fd_sc_hd__diode_2
X_0514_ _0514_/A _0810_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0846__A PAR_IN1[26] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1007__A _0809_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_234 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0581__A _0559_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0776__A1 PAR_IN3[13] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_138 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0700__A1 PAR_IN3[19] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0756__A PAR_IN5[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_142 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0666__A _0627_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_160 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_51_318 VSS VDD sky130_fd_sc_hd__fill_1
X_0994_ PAR_IN6[4] _0994_/B _0994_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0832__C _0831_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0758__A1 PAR_IN4[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_82 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_226 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_40_57 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_66 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0921__A1 _0910_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_18 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0933__B _0924_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_156 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_112 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0652__C _0652_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_80 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0912__A1 PAR_IN6[6] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_167 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_101 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1004__B _0724_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0979__A1 PAR_IN3[12] VSS VDD sky130_fd_sc_hd__diode_2
X_0977_ PAR_IN1[12] _0988_/B _0986_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_10_27 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0903__A1 PAR_IN5[22] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_159 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_27_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0737__C _0734_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0753__B _0741_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_200 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_101 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0663__B _0744_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_90 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_192 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0944__A _0944_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0900_ _0810_/A _0900_/B _0900_/C _0900_/X VSS VDD sky130_fd_sc_hd__or3_4
X_0831_ _0831_/A _0820_/X _0831_/C _0831_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_0762_ _0683_/A _0753_/X _0761_/X _0763_/C VSS VDD sky130_fd_sc_hd__and3_4
X_0693_ PAR_IN4[3] _0692_/X _0616_/X _0696_/C VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_44_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0897__B1 _0896_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_61 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0854__A _0848_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0649__B1 _0648_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1015__A _0533_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_170 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0573__B _0573_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0764__A PAR_IN1[29] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_148 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_28 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_303 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0658__B _0610_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_70 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_81 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_295 VSS VDD sky130_fd_sc_hd__fill_1
X_0814_ PAR_IN6[1] _0662_/A _0814_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0745_ PAR_IN7[5] _0645_/X _0744_/X _0745_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0567__C1 _0524_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_CLK_A CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0849__A PAR_IN6[26] VSS VDD sky130_fd_sc_hd__diode_2
X_0676_ _0656_/A _0676_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0582__A2 _0536_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_210 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0584__A _0510_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_195 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0558__C1 _0535_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0759__A PAR_IN6[21] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0909__D _0908_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_295 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_254 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0564__A2 _0561_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_184 VSS VDD sky130_fd_sc_hd__fill_2
X_0530_ _0603_/B _0524_/Y _0559_/A _0530_/D _0530_/X VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__0819__D _0818_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0669__A _0619_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_276 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_210 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1012__B COUNT[5] VSS VDD sky130_fd_sc_hd__diode_2
X_1013_ _0835_/X _1012_/X _1013_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_19_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_71 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_8_93 VSS VDD sky130_fd_sc_hd__fill_2
X_0659_ PAR_IN8[7] _0657_/X _0658_/X _0659_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0728_ PAR_IN5[11] _0694_/B _0728_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0555__A2 _0530_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_24 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_246 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_235 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0761__B _0757_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_114 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0546__A2 _0573_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_276 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_293 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_279 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_271 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0671__B _0671_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0513_ COUNT[3] _0514_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__0846__B _0591_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1007__B _1007_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0862__A PAR_IN6[18] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0581__B _0581_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0776__A2 _0725_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_68 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0700__A2 _0635_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0756__B _0749_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0772__A _0766_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_154 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_132 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0666__B _0666_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_172 VSS VDD sky130_fd_sc_hd__decap_12
X_0993_ PAR_IN4[4] _0730_/X _0732_/X _0996_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0682__A _0682_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0758__A2 _0731_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0857__A _0591_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_94 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_176 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0592__A _0924_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_205 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_102 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0921__A2 _0920_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0767__A PAR_IN5[29] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0933__C _0933_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1028__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0912__A2 _0662_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_275 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_286 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0677__A _0676_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_127 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0979__A2 _0724_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_190 VSS VDD sky130_fd_sc_hd__fill_2
X_0976_ _0976_/A _0967_/X _0976_/C _0976_/X VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_10_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0903__A2 _0789_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0737__D _0736_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_15 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0587__A SAMPLE_COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_47 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_35 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0944__B _0933_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_91 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_182 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_80 VSS VDD sky130_fd_sc_hd__decap_3
X_0830_ _0809_/A _0821_/X _0829_/X _0831_/C VSS VDD sky130_fd_sc_hd__and3_4
X_0692_ _0787_/B _0692_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0761_ _0761_/A _0757_/X _0758_/X _0761_/D _0761_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_49_271 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0897__A1 PAR_IN2[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_84 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_40 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0649__A1 PAR_IN7[31] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1015__B _1014_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0854__B _0854_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_105 VSS VDD sky130_fd_sc_hd__decap_8
X_0959_ PAR_IN8[8] _0676_/X _0958_/X _0959_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0870__A PAR_IN4[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_46 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0764__B _0741_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_108 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0780__A PAR_IN5[13] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_127 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0576__B1 _0575_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_285 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0955__A PAR_IN1[8] VSS VDD sky130_fd_sc_hd__diode_2
X_0813_ PAR_IN3[1] _0614_/X _0812_/X _0819_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0690__A PAR_IN6[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_160 VSS VDD sky130_fd_sc_hd__fill_2
X_0744_ PAR_IN6[5] _0744_/B _0744_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0675_ PAR_IN4[23] _0642_/X _0643_/X _0675_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0567__B1 _0566_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0849__B _0595_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_263 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0865__A PAR_IN8[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_37 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_141 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0558__B1 _0557_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0759__B _0597_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_233 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_43_211 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_200 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_274 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0775__A PAR_IN2[13] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_81 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0549__B1 _0548_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0685__A _1009_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1012_ SAMPLE_COUNT[3] COUNT[5] COMPLETE _1011_/Y _1012_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_19_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_230 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_34_233 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1012__C COMPLETE VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_285 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0788__B1 _0787_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1022__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
X_0727_ PAR_IN3[11] _0725_/X _0726_/X _0737_/A VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_8_83 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0960__B1 _0732_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0658_ PAR_IN5[7] _0610_/B _0658_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0589_ _0615_/A _0590_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_27_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_26 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_15 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0595__A _0595_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0779__B1 _0733_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0761__C _0758_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_19 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0703__B1 _0643_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_258 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_214 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_261 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_92 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_294 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ _0933_/A _0512_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_3_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1007__C _1007_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0862__B _0862_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_291 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0581__C READY VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0772__B _0768_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_214 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_291 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_188 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_166 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0963__A _0957_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0666__C _0665_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_195 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0682__B _0674_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0992_ PAR_IN8[4] _0676_/X _0991_/X _0992_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_5_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_133 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_111 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0915__B1 _0792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_15 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_35 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0906__B1 _0590_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_7 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0767__B _0749_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0783__A _0512_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_180 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_298 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0958__A PAR_IN5[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_90 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_125 VSS VDD sky130_fd_sc_hd__decap_8
X_0975_ _0969_/X _0971_/X _0975_/C _0974_/X _0976_/C VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0868__A COUNT[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0587__B _0587_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_224 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0944__C _0943_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_117 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_106 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_114 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_92 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_81 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_70 VSS VDD sky130_fd_sc_hd__decap_3
X_0760_ PAR_IN7[21] _0706_/X _0759_/X _0761_/D VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_41_91 VSS VDD sky130_fd_sc_hd__fill_2
X_0691_ PAR_IN7[3] _0689_/X _0690_/X _0691_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_49_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_250 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0897__A2 _0925_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0649__A2 _0645_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0854__C _0851_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_139 VSS VDD sky130_fd_sc_hd__fill_2
X_0958_ PAR_IN5[8] _0803_/B _0958_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_21_39 VSS VDD sky130_fd_sc_hd__fill_1
X_0889_ COUNT[4] _0889_/B _0889_/C _0900_/B VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0870__B _0870_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0598__A _0603_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_58 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1018__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_106 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0780__B _0749_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0576__A1 _0559_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0955__B _0988_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_264 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_172 VSS VDD sky130_fd_sc_hd__decap_8
X_0812_ PAR_IN2[1] _0956_/B _0812_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0567__A1 _1009_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0743_ PAR_IN3[5] _0725_/X _0742_/X _0751_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0690__B _0673_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_194 VSS VDD sky130_fd_sc_hd__fill_2
X_0674_ PAR_IN7[23] _0645_/X _0673_/X _0674_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_37_275 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0865__B _0852_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_131 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0881__A PAR_IN4[30] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0558__A1 _0559_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0775__B _0620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_289 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_113 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_146 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_157 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0549__A1 _0530_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_142 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_153 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_197 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0966__A COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
X_1011_ COUNT[0] _0923_/X _1010_/X _1011_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0685__B _0652_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0788__A1 PAR_IN6[9] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1012__D _1011_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0726_ PAR_IN2[11] _0671_/B _0726_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_6_190 VSS VDD sky130_fd_sc_hd__fill_2
X_0657_ _0657_/A _0657_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0960__A1 PAR_IN4[8] VSS VDD sky130_fd_sc_hd__diode_2
X_0588_ _0588_/A _0615_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_40_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_204 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0779__A1 PAR_IN4[13] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0761__D _0761_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_311 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0786__A PAR_IN1[9] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0703__A1 PAR_IN4[19] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_295 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_70 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_284 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_0511_ _0510_/X _0933_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_39_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_3_193 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0696__A _0688_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_248 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_237 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_226 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0581__D _0581_/D VSS VDD sky130_fd_sc_hd__diode_2
X_0709_ _0700_/X _0709_/B _0703_/X _0708_/X _0709_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_45_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_38_37 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_15 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0772__C _0772_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_259 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0688__B1 _0687_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_178 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0963__B _0959_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0682__C _0675_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0991_ PAR_IN5[4] _0930_/B _0991_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0915__A1 PAR_IN3[6] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_52 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0851__B1 _0615_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_49 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0906__A1 PAR_IN3[22] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0783__B _0783_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_307 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_72 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0958__B _0803_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_118 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1020__D _1020_/D VSS VDD sky130_fd_sc_hd__diode_2
X_0974_ PAR_IN8[28] _0676_/X _0973_/X _0974_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_10_19 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1010__B1 _0517_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0868__B _0868_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_28 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_39 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_310 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0794__A PAR_IN7[9] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_140 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_82 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0815__B1 _0814_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_71 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_129 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_60 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_170 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_71 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_126 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_184 VSS VDD sky130_fd_sc_hd__fill_2
X_0690_ PAR_IN6[3] _0673_/B _0690_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1016__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_97 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_53 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0854__D _0853_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_140 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_192 VSS VDD sky130_fd_sc_hd__fill_1
X_0957_ PAR_IN3[8] _0614_/X _0956_/X _0957_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0879__A _0944_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0888_ _0888_/A _0888_/B _0888_/C _0887_/X _0889_/C VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0598__B SAMPLE_COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0576__A2 _0573_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_84 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0789__A _0608_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_151 VSS VDD sky130_fd_sc_hd__fill_2
X_0673_ PAR_IN6[23] _0673_/B _0673_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_52_80 VSS VDD sky130_fd_sc_hd__fill_2
X_0811_ PAR_IN1[1] _0988_/B _0811_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0567__A2 _0519_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0699__A PAR_IN2[19] VSS VDD sky130_fd_sc_hd__diode_2
X_0742_ PAR_IN2[5] _0671_/B _0742_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_42_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_224 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_20_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0881__B _0870_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0558__A2 COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_290 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_110 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0549__A2 _0547_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_176 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0966__B _0944_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_91 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_257 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_224 VSS VDD sky130_fd_sc_hd__decap_3
X_1010_ _0966_/Y _1009_/Y _0517_/Y _1010_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__0685__C _0684_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0788__A2 _0744_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0960__A2 _0692_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0725_ _0724_/X _0725_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0656_ _0656_/A _0657_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_27_39 VSS VDD sky130_fd_sc_hd__fill_2
X_0587_ SAMPLE_COUNT[3] _0587_/B _0588_/A VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_43_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_235 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0779__A2 _0731_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_316 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0786__B _0967_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0703__A2 _0642_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_213 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_296 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_82 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_274 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_0510_ _0509_/Y _0510_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_3_150 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0977__A PAR_IN1[12] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0696__B _0691_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1023__D _1023_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_19 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_27 VSS VDD sky130_fd_sc_hd__decap_4
X_0708_ PAR_IN7[19] _0706_/X _0707_/X _0708_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0639_ PAR_IN3[31] _0635_/X _0638_/X _0639_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_38_49 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_9_209 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0772__D _0771_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_249 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_102 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0797__A _0933_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0688__A1 PAR_IN3[3] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0963__C _0963_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0682__D _0682_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_93 VSS VDD sky130_fd_sc_hd__fill_2
X_0990_ PAR_IN3[4] _0724_/X _0989_/X _0990_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_8_242 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_260 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0915__A2 _0724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_97 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1018__D _0581_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_157 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_146 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0851__A1 PAR_IN3[26] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0906__A2 _0724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0783__C _0783_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_84 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_83 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_182 VSS VDD sky130_fd_sc_hd__fill_2
X_0973_ PAR_IN5[28] _0803_/B _0973_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1010__A1 _0966_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0868__C _0867_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_108 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_171 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_149 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_300 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_27 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_204 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0794__B _0794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_138 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0760__B1 _0759_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_94 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_83 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_163 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0815__A1 PAR_IN7[1] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_72 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_61 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_182 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_50 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_196 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_71 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0579__B1 _0578_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0985__A _0985_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_32 VSS VDD sky130_fd_sc_hd__decap_8
X_0956_ PAR_IN2[8] _0956_/B _0956_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_32_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_130 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_19 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0990__B1 _0989_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0887_ PAR_IN2[30] _0925_/B _0886_/X _0887_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0879__B _0879_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0598__C _0603_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_130 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0981__B1 _0980_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_11_74 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_71 VSS VDD sky130_fd_sc_hd__decap_12
X_0810_ _0810_/A _0810_/B _0809_/X _0810_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_36_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0972__B1 _0792_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0699__B _0699_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0741_ PAR_IN1[5] _0741_/B _0741_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0672_ PAR_IN3[23] _0635_/X _0671_/X _0682_/A VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_37_233 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1026__D _0549_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_258 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_236 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_19 VSS VDD sky130_fd_sc_hd__fill_2
X_0939_ PAR_IN4[16] _0600_/X _0792_/X _0939_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_32_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_177 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_166 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_299 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_244 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_233 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_40 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_310 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0966__C _0965_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_233 VSS VDD sky130_fd_sc_hd__fill_2
X_0724_ _0724_/A _0724_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0655_ PAR_IN3[7] _0635_/X _0654_/X _0665_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0586_ _0586_/A _0586_/B _0618_/B _0587_/B VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_25_214 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_269 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_225 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0936__B1 _0935_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_206 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_247 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_73 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_297 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0977__B _0988_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_173 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0696__C _0696_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0707_ PAR_IN6[19] _0744_/B _0707_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0569_ _0559_/X _0567_/X _0568_/X _1021_/D VSS VDD sky130_fd_sc_hd__a21oi_4
X_0638_ PAR_IN2[31] _0699_/B _0638_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0797__B _0786_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_136 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_83 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_61 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0688__A2 _0614_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_187 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_93 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0963__D _0962_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_221 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_276 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_298 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0988__A PAR_IN1[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_103 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_169 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0851__A2 _0842_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_19 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0898__A _0898_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_49 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_224 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_60 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0601__A PAR_IN4[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_194 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_172 VSS VDD sky130_fd_sc_hd__fill_2
X_0972_ PAR_IN4[28] _0600_/X _0792_/X _0975_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0511__A _0510_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1010__A2 _1009_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_290 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_150 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_39 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_164 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_249 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0760__A1 PAR_IN7[21] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_95 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_84 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_131 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0815__A2 _0705_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_73 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_62 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_51 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_95 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_25_62 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_40 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_9 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0579__A1 _0559_/X VSS VDD sky130_fd_sc_hd__diode_2
Xclkbuf_0_CLK CLK clkbuf_0_CLK/X VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_49_275 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0985__B _0985_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_282 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_297 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_161 VSS VDD sky130_fd_sc_hd__decap_3
X_0955_ PAR_IN1[8] _0988_/B _0955_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0886_ PAR_IN8[30] _0852_/B _0886_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1025__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0990__A1 PAR_IN3[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0879__C _0879_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0598__D _0618_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0981__A1 PAR_IN8[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_234 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_83 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_131 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_93 VSS VDD sky130_fd_sc_hd__fill_2
X_0740_ COUNT[2] _0740_/B _0740_/C _0740_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_14_164 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0996__A _0990_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0972__A1 PAR_IN4[28] VSS VDD sky130_fd_sc_hd__diode_2
X_0671_ PAR_IN2[23] _0671_/B _0671_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_37_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0660__B1 _0643_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0869_ PAR_IN1[2] _0901_/B _0869_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0938_ PAR_IN8[16] _0657_/A _0937_/X _0938_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_28_289 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_189 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_71 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_245 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_201 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_237 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_289 VSS VDD sky130_fd_sc_hd__decap_12
X_0723_ PAR_IN1[11] _0741_/B _0723_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_8_32 VSS VDD sky130_fd_sc_hd__fill_2
X_0654_ PAR_IN2[7] _0699_/B _0654_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0585_ SAMPLE_COUNT[2] _0618_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_25_259 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0936__A1 PAR_IN3[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_218 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_243 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_281 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_232 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_85 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_298 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_276 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0604__A _0852_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0696__D _0695_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0863__B1 _0862_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0514__A _0514_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0706_ _0705_/X _0706_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0568_ _0550_/X _1009_/A _0562_/X _0568_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0637_ _0637_/A _0699_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_13_207 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_218 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0797__C _0796_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_72 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_8_211 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0988__B _0988_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_137 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_115 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0509__A COUNT[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0898__B _0898_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_195 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_203 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_5_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_258 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0601__B _0600_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0818__B1 _0817_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_107 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_302 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_17_310 VSS VDD sky130_fd_sc_hd__decap_8
X_0971_ PAR_IN7[28] _0645_/A _0970_/X _0971_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0999__A PAR_IN7[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_154 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_198 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_176 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0760__A2 _0706_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_228 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_129 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_30 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_96 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_85 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_74 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_63 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0579__A2 _0524_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_52 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_41 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_41 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_95 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0612__A _0618_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_221 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0985__C _0982_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_165 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_195 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_184 VSS VDD sky130_fd_sc_hd__decap_8
X_0954_ _0976_/A _0945_/X _0953_/X _0954_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0885_ PAR_IN3[30] _0634_/A _0590_/A _0888_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0990__A2 _0724_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0981__A2 _0657_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0607__A _0618_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_72 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_61 VSS VDD sky130_fd_sc_hd__fill_1
X_0670_ _0946_/B _0671_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_14_198 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0996__B _0992_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0972__A2 _0600_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_279 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_37_213 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0660__A1 PAR_IN4[7] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0517__A COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
X_0799_ PAR_IN1[25] _0988_/B _0799_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0868_ COUNT[4] _0868_/B _0867_/X _0879_/B VSS VDD sky130_fd_sc_hd__and3_4
X_0937_ PAR_IN5[16] _0930_/B _0937_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_43_205 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_268 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_271 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_3_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_257 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_224 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_213 VSS VDD sky130_fd_sc_hd__decap_4
X_0653_ PAR_IN1[7] _0631_/X _0666_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_6_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_172 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_194 VSS VDD sky130_fd_sc_hd__decap_12
X_0722_ _0593_/B _0741_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0584_ _0510_/X _0627_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_40_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0800__A _0619_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_208 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_25_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_205 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_219 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0936__A2 _0634_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0710__A _0683_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_304 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_308 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_277 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0620__A _0925_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0560__B1 _0519_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_197 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_131 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0863__A1 PAR_IN7[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_274 VSS VDD sky130_fd_sc_hd__fill_1
X_0705_ _0794_/B _0705_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1021__CLK _1022_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_0636_ _0619_/A _0637_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0530__A _0603_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0567_ _1009_/A _0519_/B _0566_/Y _0524_/Y _0567_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_53_311 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0705__A _0794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_52 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_84 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_51 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0615__A _0615_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_234 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_245 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_296 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0781__B1 _0780_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_56 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_193 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1019__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0525__A SAMPLE_COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
X_0619_ _0619_/A _0925_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0898__C _0898_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_76 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_86 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_39_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_141 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0818__A1 PAR_IN8[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_314 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_171 VSS VDD sky130_fd_sc_hd__fill_2
X_0970_ PAR_IN6[28] _0646_/X _0970_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0999__B _0794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_133 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_122 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_196 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_314 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0993__B1 _0732_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0745__B1 _0744_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_64 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_53 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_53 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_42 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_20 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_31 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_97 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0984__B1 _0983_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_86 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_155 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_52 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_30 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_75 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_75 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0736__B1 _0735_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0612__B _0618_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_266 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_233 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0985__D _0984_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_68 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_152 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0803__A PAR_IN5[25] VSS VDD sky130_fd_sc_hd__diode_2
X_0953_ _0953_/A _0953_/B _0950_/X _0953_/D _0953_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0884_ PAR_IN7[30] _0794_/B _0883_/X _0888_/B VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0727__B1 _0726_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_155 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0713__A PAR_IN2[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_77 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_99 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_40 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0607__B _0581_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_84 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0957__B1 _0956_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0623__A _0623_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0996__C _0996_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_206 VSS VDD sky130_fd_sc_hd__fill_2
X_0936_ PAR_IN3[16] _0634_/X _0935_/X _0936_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0660__A2 _0642_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_158 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_103 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0533__A _0533_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0798_ _0924_/B _0988_/B VSS VDD sky130_fd_sc_hd__buf_1
X_0867_ _0867_/A _0863_/X _0864_/X _0866_/X _0867_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_28_236 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_258 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_103 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_294 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0939__B1 _0792_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_98 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_87 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_32 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_95 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0618__A _0618_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_67 VSS VDD sky130_fd_sc_hd__fill_2
X_0652_ _0965_/A _0627_/X _0652_/C _0652_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_6_162 VSS VDD sky130_fd_sc_hd__decap_4
X_0721_ _0683_/A _0721_/B _0721_/C _0739_/B VSS VDD sky130_fd_sc_hd__and3_4
X_0583_ _0534_/X _0583_/B _1017_/D VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_33_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_280 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0528__A COMPLETE VSS VDD sky130_fd_sc_hd__diode_2
X_0919_ PAR_IN1[6] _0924_/B _0509_/Y _0919_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_33_283 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0710__B _0710_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_54 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_289 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_278 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_53 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_267 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0901__A PAR_IN1[22] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0560__A1 COUNT[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_8 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0863__A2 _0623_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_283 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0811__A PAR_IN1[1] VSS VDD sky130_fd_sc_hd__diode_2
X_0566_ _0519_/X _0566_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_0635_ _0634_/X _0635_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0704_ _0896_/B _0794_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0530__B _0524_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_297 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0721__A _0683_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_106 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_97 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_86 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_75 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_264 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0631__A _0967_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0781__A1 PAR_IN8[13] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0806__A PAR_IN6[25] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0541__A SAMPLE_COUNT[3] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0898__D _0897_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0618_ _0618_/A _0618_/B _0618_/C _0603_/B _0619_/A VSS VDD sky130_fd_sc_hd__and4_4
X_0549_ _0530_/D _0547_/X _0548_/X _0549_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_38_194 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_183 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_38_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_52 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_150 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_186 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0626__A _0626_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0818__A2 _0606_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_101 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_175 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0536__A _0559_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0745__A1 PAR_IN7[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 PAR_IN4[4] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_98 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_87 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_123 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_76 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_65 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0681__B1 _0680_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_54 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_87 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_43 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_10 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_32 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0984__A1 PAR_IN7[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_75 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0612__C _0603_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0736__A1 PAR_IN7[11] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_263 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_131 VSS VDD sky130_fd_sc_hd__fill_1
X_0952_ PAR_IN8[24] _0606_/X _0951_/X _0953_/D VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_32_189 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0672__B1 _0671_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_175 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0803__B _0803_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0727__A1 PAR_IN3[11] VSS VDD sky130_fd_sc_hd__diode_2
X_0883_ PAR_IN6[30] _0862_/B _0883_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_23_145 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_112 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0713__B _0671_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_248 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_215 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0904__A PAR_IN6[22] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0607__C _0618_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_112 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_134 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0957__A1 PAR_IN3[8] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0996__D _0995_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_8 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_259 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0814__A PAR_IN6[1] VSS VDD sky130_fd_sc_hd__diode_2
X_0935_ PAR_IN2[16] _0946_/B _0935_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0866_ PAR_IN2[18] _0637_/A _0865_/X _0866_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_9_182 VSS VDD sky130_fd_sc_hd__fill_1
X_0797_ _0933_/A _0786_/X _0796_/X _0810_/B VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_28_215 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_204 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0884__B1 _0883_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_229 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0724__A _0724_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0939__A1 PAR_IN4[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_11 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_85 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_237 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0618__B _0618_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0634__A _0634_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0720_ _0714_/X _0720_/B _0717_/X _0719_/X _0721_/C VSS VDD sky130_fd_sc_hd__or4_4
X_0651_ _0809_/A _0651_/B _0650_/X _0652_/C VSS VDD sky130_fd_sc_hd__and3_4
X_0582_ _0535_/X _0536_/X _0530_/D _0531_/Y _0583_/B VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__0809__A _0809_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_3 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0866__B1 _0865_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_229 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_25_218 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_270 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0544__A SAMPLE_COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
X_0918_ _0912_/X _0914_/X _0915_/X _0918_/D _0918_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0849_ PAR_IN6[26] _0595_/A _0849_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0710__C _0709_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_207 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_77 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_279 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_295 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_235 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0901__B _0901_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0629__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0848__B1 _0847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0560__A2 COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_221 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0811__B _0988_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_276 VSS VDD sky130_fd_sc_hd__fill_2
X_0703_ PAR_IN4[19] _0642_/X _0643_/X _0703_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0565_ _0515_/Y _1009_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0634_ _0634_/A _0634_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0530__C _0559_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_210 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0721__B _0721_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_118 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_29_310 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_125 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_64 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_225 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_12_232 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_276 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0781__A2 _0677_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_316 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0806__B _0994_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1028__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0822__A PAR_IN2[17] VSS VDD sky130_fd_sc_hd__diode_2
X_0617_ PAR_IN3[15] _0614_/X _0616_/X _0617_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0548_ _0618_/C _0535_/X _0534_/X _0548_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_53_198 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_187 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0732__A _0792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_11 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_23 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_31 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_66 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_86 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_75 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0907__A PAR_IN8[22] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_198 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_44_176 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0626__B _0611_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0642__A _0600_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_154 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_132 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0817__A PAR_IN5[1] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0536__B _0573_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_168 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0993__A2 _0730_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0552__A _0552_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0745__A2 _0645_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_99 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_88 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_113 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_77 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_66 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_55 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0681__A1 PAR_IN8[23] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_33 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_11 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_44 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_11 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_33 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0984__A2 _0705_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_87 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0612__D _0621_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_224 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0736__A2 _0706_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_15 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_286 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_1_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_220 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_279 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_102 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0637__A _0637_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_143 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_121 VSS VDD sky130_fd_sc_hd__fill_1
X_0951_ PAR_IN5[24] _0803_/B _0951_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_40_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0672__A1 PAR_IN3[23] VSS VDD sky130_fd_sc_hd__diode_2
X_0882_ PAR_IN5[30] _0789_/X _0881_/X _0888_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0727__A2 _0725_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0547__A _0577_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_35 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_205 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_32 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_20 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0957__A2 _0614_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_190 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0904__B _0862_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0607__D _0621_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_282 VSS VDD sky130_fd_sc_hd__decap_4
X_0934_ PAR_IN1[16] _0967_/B _0934_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0814__B _0662_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_127 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0830__A _0809_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0865_ PAR_IN8[18] _0852_/B _0865_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0796_ _0788_/X _0791_/X _0796_/C _0795_/X _0796_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1024__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_227 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0884__A1 PAR_IN7[30] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_285 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_263 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_127 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_138 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_149 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0939__A2 _0600_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_45 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0740__A COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_42 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0572__B1 _0520_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_205 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_47_75 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_263 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_230 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0618__C _0618_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0650__A _0639_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_36 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_182 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_193 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0563__B1 _0562_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0581_ _0559_/X _0581_/B READY _0581_/D _0581_/X VSS VDD sky130_fd_sc_hd__and4_4
X_0650_ _0639_/X _0650_/B _0644_/X _0649_/X _0650_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_6_186 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0809__B _0799_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0866__A1 PAR_IN2[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_241 VSS VDD sky130_fd_sc_hd__decap_3
X_0848_ PAR_IN5[26] _0747_/A _0847_/X _0848_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0917_ PAR_IN2[6] _0699_/B _0916_/X _0918_/D VSS VDD sky130_fd_sc_hd__a21o_4
X_0779_ PAR_IN4[13] _0731_/X _0733_/X _0779_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_24_252 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0735__A PAR_IN6[11] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_225 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_66 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_269 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_236 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0793__B1 _0792_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_300 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0848__A1 PAR_IN5[26] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0645__A _0645_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_233 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_263 VSS VDD sky130_fd_sc_hd__decap_12
X_0702_ PAR_IN8[19] _0657_/X _0701_/X _0709_/B VSS VDD sky130_fd_sc_hd__a21o_4
X_0633_ _0842_/B _0634_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0564_ _0559_/X _0561_/Y _0563_/X _1020_/D VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__0530__D _0530_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_81 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_222 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0721__C _0721_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_137 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0766__B1 _0765_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_48 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_163 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0822__B _0956_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0616_ _0792_/A _0616_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0757__B1 _0756_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0547_ _0577_/A _0547_/B _0547_/C _0547_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_41_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_68 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_133 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0907__B _0907_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0920__B1 _0944_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_196 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0626__C _0617_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0923__A COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_251 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0817__B _0610_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0833__A COUNT[1] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0552__B _0547_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_133 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_12 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_89 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0969__B1 _0968_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_136 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_78 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_67 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_56 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0681__A2 _0677_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_56 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_45 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_23 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_306 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_34 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_99 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_258 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0918__A _0912_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_298 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_254 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0672__A2 _0635_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_166 VSS VDD sky130_fd_sc_hd__fill_2
X_0950_ PAR_IN4[24] _0730_/X _0792_/X _0950_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_32_158 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0653__A PAR_IN1[7] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_309 VSS VDD sky130_fd_sc_hd__decap_8
X_0881_ PAR_IN4[30] _0870_/B _0881_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_49_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_291 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0547__B _0547_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_191 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0738__A _0512_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_43 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_32 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0648__A PAR_IN6[31] VSS VDD sky130_fd_sc_hd__diode_2
X_0933_ _0933_/A _0924_/X _0933_/C _0933_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0795_ PAR_IN2[9] _0620_/X _0794_/X _0795_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0864_ PAR_IN3[18] _0634_/A _0615_/A _0864_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_9_184 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0830__B _0821_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_92 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_272 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0884__A2 _0794_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0572__A1 _0831_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0740__B _0740_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_21 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_217 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_261 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0618__D _0603_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0650__B _0650_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_90 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0563__A1 _0550_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0580_ _0550_/X _0530_/D COUNT[5] _0533_/A _0580_/X VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__0809__C _0809_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0866__A2 _0637_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_250 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_275 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_253 VSS VDD sky130_fd_sc_hd__fill_2
X_0916_ PAR_IN7[6] _0623_/A _0916_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0847_ PAR_IN4[26] _0599_/A _0847_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0778_ PAR_IN7[13] _0706_/X _0777_/X _0778_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_33_34 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_259 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0735__B _0744_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_226 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_68 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0793__A1 PAR_IN3[9] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_89 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0751__A _0751_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_113 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0848__A2 _0747_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0661__A _0862_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_275 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_297 VSS VDD sky130_fd_sc_hd__fill_2
X_0563_ _0550_/X _0517_/Y _0562_/X _0563_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0632_ PAR_IN1[31] _0631_/X _0651_/B VSS VDD sky130_fd_sc_hd__or2_4
X_0701_ PAR_IN5[19] _0694_/B _0701_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_31_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_53_304 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0836__A PAR_IN1[10] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0571__A _0944_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_267 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_80 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_0_149 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_56 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_256 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_27 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_38 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0766__A1 PAR_IN3[29] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0656__A _0656_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0757__A1 PAR_IN8[21] VSS VDD sky130_fd_sc_hd__diode_2
X_0615_ _0615_/A _0792_/A VSS VDD sky130_fd_sc_hd__buf_1
X_0546_ _0621_/D _0573_/A _0618_/C _0547_/C VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_38_186 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_142 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_131 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_120 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0566__A _0519_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_156 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_36 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0693__B1 _0616_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_79 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_11 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0920__A1 _0918_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_112 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0626__D _0625_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_29_175 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0923__B _0922_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_230 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_137 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0675__B1 _0643_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0833__B _0832_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_318 VSS VDD sky130_fd_sc_hd__fill_1
X_0529_ _0552_/A _0530_/D VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_26_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_112 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_46 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_35 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_13 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0969__A1 PAR_IN3[28] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_159 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_56 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_79 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_68 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_57 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_68 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_237 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0918__B _0914_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0934__A PAR_IN1[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_148 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0653__B _0631_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_123 VSS VDD sky130_fd_sc_hd__decap_8
X_0880_ PAR_IN1[30] _0901_/B _0889_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_23_104 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0547__C _0547_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0844__A _0838_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_159 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_270 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0887__B1 _0886_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0738__B _0723_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_292 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_45 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0754__A PAR_IN2[21] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0639__B1 _0638_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_303 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0648__B _0673_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0932_ _0932_/A _0928_/X _0929_/X _0931_/X _0933_/C VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_20_118 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0802__B1 _0801_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0794_ PAR_IN7[9] _0794_/B _0794_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0863_ PAR_IN7[18] _0623_/A _0862_/X _0863_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0830__C _0829_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_163 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_196 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0839__A PAR_IN6[10] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0574__A _0810_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_262 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_118 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0749__A PAR_IN5[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0572__A2 _0566_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0740__C _0740_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_99 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_47_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_287 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_243 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_27 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0650__C _0644_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_8 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0563__A2 _0517_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_284 VSS VDD sky130_fd_sc_hd__decap_12
X_0915_ PAR_IN3[6] _0724_/A _0792_/A _0915_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0846_ PAR_IN1[26] _0591_/A _0846_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0777_ PAR_IN6[13] _0597_/X _0777_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_17_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_57 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_249 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_287 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_24_276 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_227 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_58 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0793__A2 _0724_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0751__B _0745_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_169 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_232 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0942__A _0936_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_246 VSS VDD sky130_fd_sc_hd__decap_12
X_0700_ PAR_IN3[19] _0635_/X _0699_/X _0700_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0631_ _0967_/B _0631_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0562_ COMPLETE _0562_/B _0562_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_24_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0836__B _0591_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0852__A PAR_IN8[26] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1013__A _0835_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_94 VSS VDD sky130_fd_sc_hd__decap_12
X_0829_ _0823_/X _0829_/B _0826_/X _0829_/D _0829_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_0_106 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_79 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_46 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0762__A _0683_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_202 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_290 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0766__A2 _0725_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_132 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0937__A PAR_IN5[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_308 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0757__A2 _0677_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1008__A _0944_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0614_ _0724_/A _0614_/X VSS VDD sky130_fd_sc_hd__buf_1
X_0545_ _0586_/A _0618_/C VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0847__A PAR_IN4[26] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_198 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_154 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0693__A1 PAR_IN4[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_168 VSS VDD sky130_fd_sc_hd__decap_12
X_1028_ _0556_/X SAMPLE_COUNT[3] RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_14_26 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_47 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_34 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0920__A2 _0919_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_168 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0675__A1 PAR_IN4[23] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0667__A _0809_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_149 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_105 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_157 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1027__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0577__A _0577_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0528_ COMPLETE _0552_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_41_127 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_69 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_14 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_47 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_36 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_14 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0969__A2 _0634_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_79 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_41_24 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_13 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0918__C _0915_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_113 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_278 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0934__B _0967_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_179 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_157 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_80 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_48_271 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0844__B _0840_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_171 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_160 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0860__A PAR_IN4[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_13 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1021__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0887__A1 PAR_IN2[30] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0738__C _0737_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0639__A1 PAR_IN3[31] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0754__B _0671_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_127 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0770__A PAR_IN6[29] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_182 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_315 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0575__B1 _0562_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0945__A PAR_IN1[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_219 VSS VDD sky130_fd_sc_hd__fill_2
X_0931_ PAR_IN8[0] _0657_/A _0930_/X _0931_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0680__A PAR_IN5[23] VSS VDD sky130_fd_sc_hd__diode_2
X_0862_ PAR_IN6[18] _0862_/B _0862_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0802__A1 PAR_IN3[25] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_193 VSS VDD sky130_fd_sc_hd__fill_2
X_0793_ PAR_IN3[9] _0724_/X _0792_/X _0796_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0839__B _0595_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_222 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0855__A COUNT[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_241 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0590__A _0590_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0749__B _0749_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0557__B1 _0518_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_67 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_208 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0765__A PAR_IN2[29] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_299 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_10_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0650__D _0649_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0548__B1 _0534_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_296 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_263 VSS VDD sky130_fd_sc_hd__decap_4
X_0845_ _0510_/X _0836_/X _0844_/X _0845_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0914_ PAR_IN8[6] _0656_/A _0913_/X _0914_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0776_ PAR_IN3[13] _0725_/X _0775_/X _0782_/A VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0539__B1 _0621_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0585__A SAMPLE_COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_239 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_299 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_244 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0751__C _0751_/C VSS VDD sky130_fd_sc_hd__diode_2
XPHY_228 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0778__B1 _0777_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0950__B1 _0792_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0702__B1 _0701_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_200 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0942__B _0938_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_258 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_30_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_91 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0769__B1 _0733_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_288 VSS VDD sky130_fd_sc_hd__fill_2
X_0630_ _0924_/B _0967_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0941__B1 _0940_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0561_ _0573_/A _0560_/X _0561_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_0_40 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0852__B _0852_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1013__B _1012_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_236 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_214 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_203 VSS VDD sky130_fd_sc_hd__decap_4
X_0759_ PAR_IN6[21] _0597_/X _0759_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0828_ PAR_IN7[17] _0689_/X _0827_/X _0829_/D VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_29_314 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_118 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_13 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0762__B _0753_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_229 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_306 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0937__B _0930_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0953__A _0953_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0613_ _0842_/B _0724_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_295 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0847__B _0599_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1008__B _0997_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0914__B1 _0913_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0544_ SAMPLE_COUNT[1] _0586_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_53_125 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_177 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_166 VSS VDD sky130_fd_sc_hd__fill_2
X_1027_ _0555_/Y SAMPLE_COUNT[2] RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0693__A2 _0692_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0905__B1 _0904_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_188 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0773__A _0683_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0948__A PAR_IN6[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_298 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_114 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0675__A2 _0642_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0683__A _0683_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_117 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0577__B _0520_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0858__A PAR_IN1[18] VSS VDD sky130_fd_sc_hd__diode_2
X_0527_ _0618_/A _0559_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0593__A PAR_IN1[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_117 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_59 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_158 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_37 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_48 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_37 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_217 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_224 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0918__D _0918_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_103 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_106 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0678__A _0747_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0844__C _0844_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_150 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0860__B _0870_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0588__A _0588_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0887__A2 _0925_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0639__A2 _0635_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_68 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_194 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_139 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0770__B _0597_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0575__A1 _0577_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_264 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0945__B _0967_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1017__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_0930_ PAR_IN5[0] _0930_/B _0930_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0802__A2 _0724_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0680__B _0694_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0961__A PAR_IN6[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_90 VSS VDD sky130_fd_sc_hd__fill_2
X_0792_ _0792_/A _0792_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_20_109 VSS VDD sky130_fd_sc_hd__fill_2
X_0861_ PAR_IN5[18] _0789_/X _0860_/X _0867_/A VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_9_132 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_40 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0855__B _0846_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0557__A1 _0577_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_201 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_297 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_264 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_253 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0765__B _0620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_267 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_102 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_124 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_186 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_146 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_168 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0548__A1 _0618_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0956__A PAR_IN2[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_7 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_234 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_201 VSS VDD sky130_fd_sc_hd__fill_2
X_0844_ _0838_/X _0840_/X _0844_/C _0844_/D _0844_/X VSS VDD sky130_fd_sc_hd__or4_4
X_0913_ PAR_IN5[6] _0747_/A _0913_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0775_ PAR_IN2[13] _0620_/X _0775_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0539__A1 _0535_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_201 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_207 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_49 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0751__D _0750_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0778__A1 PAR_IN7[13] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_256 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_229 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_105 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0950__A1 PAR_IN4[24] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_304 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0702__A1 PAR_IN8[19] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0942__C _0939_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_81 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_70 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0769__A1 PAR_IN4[29] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0941__A1 PAR_IN7[16] VSS VDD sky130_fd_sc_hd__diode_2
X_0560_ COUNT[0] COUNT[1] _0519_/B _0560_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_2_182 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0686__A PAR_IN1[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_63 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_9_50 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_83 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_94 VSS VDD sky130_fd_sc_hd__fill_2
X_0758_ PAR_IN4[21] _0731_/X _0733_/X _0758_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0827_ PAR_IN6[17] _0673_/B _0827_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0689_ _0645_/A _0689_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0596__A _0862_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_44_47 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0762__C _0761_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_19 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_167 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0953__B _0953_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_91 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0611__B1 _0610_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_230 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_281 VSS VDD sky130_fd_sc_hd__fill_2
X_0612_ _0618_/A _0618_/B _0603_/A _0621_/D _0842_/B VSS VDD sky130_fd_sc_hd__and4_4
XFILLER_38_101 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1008__C _1008_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0914__A1 PAR_IN8[6] VSS VDD sky130_fd_sc_hd__diode_2
X_0543_ _0603_/A _0603_/B _0524_/Y _0547_/B VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_53_137 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_307 VSS VDD sky130_fd_sc_hd__decap_12
X_1026_ _0549_/Y SAMPLE_COUNT[1] RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0602__B1 _0601_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0850__B1 _0849_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_25 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0905__A1 PAR_IN7[22] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_137 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_69 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_101 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_44_159 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0841__B1 _0615_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0773__B _0773_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0948__B _0662_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_93 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0964__A _0627_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0683__B _0668_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0858__B _0901_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_51 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_6_73 VSS VDD sky130_fd_sc_hd__decap_12
X_0526_ _0603_/C _0618_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0593__B _0593_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1009_ _1009_/A _0987_/Y _1009_/C _1009_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_25_49 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_49 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_38 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0823__B1 _0822_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_16 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_48 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_236 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1000__B1 _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_118 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0784__A _0965_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_148 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_162 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_140 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_310 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_92 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_70 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0694__A PAR_IN5[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_280 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0805__B1 _0732_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0844__D _0844_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_195 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_29 VSS VDD sky130_fd_sc_hd__decap_4
X_0509_ COUNT[4] _0509_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__0869__A PAR_IN1[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_37 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0575__A2 _0965_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_243 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_221 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0961__B _0994_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0791_ PAR_IN8[9] _0657_/A _0790_/X _0791_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0860_ PAR_IN4[18] _0870_/B _0860_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_13_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0689__A _0645_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_202 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0855__C _0854_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_276 VSS VDD sky130_fd_sc_hd__decap_8
X_0989_ PAR_IN2[4] _0946_/B _0989_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0599__A _0599_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0557__A2 COUNT[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_235 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_232 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_114 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_136 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_158 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_110 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_61 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0548__A2 _0535_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0956__B _0956_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_276 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_210 VSS VDD sky130_fd_sc_hd__decap_4
X_0912_ PAR_IN6[6] _0662_/A _0911_/X _0912_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_33_279 VSS VDD sky130_fd_sc_hd__fill_2
X_0843_ PAR_IN5[10] _0789_/X _0842_/X _0844_/D VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0539__A2 _0536_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0774_ PAR_IN1[13] _0741_/B _0783_/B VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_24_268 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_213 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_219 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0778__A2 _0706_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0950__A2 _0730_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_117 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0702__A2 _0657_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0942__D _0941_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0792__A _0792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_290 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_279 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0769__A2 _0731_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0967__A PAR_IN1[28] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_305 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0941__A2 _0705_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0686__B _0593_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_40 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_62 VSS VDD sky130_fd_sc_hd__decap_12
X_0688_ PAR_IN3[3] _0614_/X _0687_/X _0688_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0877__A _0871_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0757_ PAR_IN8[21] _0677_/X _0756_/X _0757_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_0_109 VSS VDD sky130_fd_sc_hd__decap_3
X_0826_ PAR_IN4[17] _0692_/X _0616_/X _0826_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_44_59 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0787__A PAR_IN4[9] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_113 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0953__C _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_260 VSS VDD sky130_fd_sc_hd__fill_2
X_0611_ PAR_IN8[15] _0606_/X _0610_/X _0611_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0611__A1 PAR_IN8[15] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0914__A2 _0656_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0542_ SAMPLE_COUNT[1] _0603_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_264 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_135 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0697__A _0627_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_149 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0850__A1 PAR_IN7[26] VSS VDD sky130_fd_sc_hd__diode_2
X_1025_ _0540_/Y SAMPLE_COUNT[0] RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_0809_ _0809_/A _0799_/X _0809_/C _0809_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0602__A1 PAR_IN6[15] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0905__A2 _0794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_105 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_179 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0773__C _0773_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0841__A1 PAR_IN8[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_72 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_223 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_234 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_160 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0964__B _0955_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0980__A PAR_IN5[12] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0683__C _0683_/C VSS VDD sky130_fd_sc_hd__diode_2
XPHY_380 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VSS VDD sky130_fd_sc_hd__decap_6
X_0525_ SAMPLE_COUNT[3] _0603_/C VSS VDD sky130_fd_sc_hd__inv_8
XPHY_17 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_28 VSS VDD sky130_fd_sc_hd__decap_3
X_1008_ _0944_/A _0997_/X _1008_/C _1009_/C VSS VDD sky130_fd_sc_hd__nor3_4
XPHY_39 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0823__A1 PAR_IN3[17] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0890__A PAR_IN1[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_259 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1000__A1 PAR_IN5[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_182 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0784__B _0784_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_185 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0578__B1 _0562_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0694__B _0694_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_296 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_241 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0975__A _0969_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0750__B1 _0749_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_292 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0805__A1 PAR_IN4[25] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1021__D _1021_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_23_108 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_171 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0569__B1 _0568_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0869__B _0901_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0508_ SAMPLE_COUNT[0] _0603_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_39_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_163 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_130 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_93 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_130 VSS VDD sky130_fd_sc_hd__fill_2
X_0790_ PAR_IN5[9] _0789_/X _0790_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_9_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_178 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0971__B1 _0970_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_53 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1016__D _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_244 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_222 VSS VDD sky130_fd_sc_hd__decap_4
X_0988_ PAR_IN1[4] _0988_/B _0988_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0962__B1 _0961_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_200 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0714__B1 _0713_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_247 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_280 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_122 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_84 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_280 VSS VDD sky130_fd_sc_hd__decap_4
X_0911_ PAR_IN4[6] _0787_/B _0911_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0842_ PAR_IN3[10] _0842_/B _0842_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_52_3 VSS VDD sky130_fd_sc_hd__decap_8
X_0773_ _0683_/A _0773_/B _0773_/C _0784_/B VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_33_28 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_209 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_30_206 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0926__B1 _0925_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0967__B _0967_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_7 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_151 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0983__A PAR_IN6[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_32 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_43 VSS VDD sky130_fd_sc_hd__fill_2
X_0825_ PAR_IN8[17] _0606_/X _0824_/X _0829_/B VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_9_74 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0917__B1 _0916_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0877__B _0873_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0756_ PAR_IN5[21] _0749_/B _0756_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0687_ PAR_IN2[3] _0699_/B _0687_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_29_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_17 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0893__A PAR_IN5[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_228 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0908__B1 _0907_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_294 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0787__B _0787_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0953__D _0953_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0611__A2 _0606_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_272 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_50_81 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0978__A PAR_IN2[12] VSS VDD sky130_fd_sc_hd__diode_2
X_0610_ PAR_IN5[15] _0610_/B _0610_/X VSS VDD sky130_fd_sc_hd__and2_4
X_0541_ SAMPLE_COUNT[3] _0577_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0697__B _0697_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_106 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1024__D _0580_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1024_ _0580_/X COUNT[5] RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_15_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0850__A2 _0623_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_19 VSS VDD sky130_fd_sc_hd__decap_4
X_0808_ _0808_/A _0804_/X _0805_/X _0807_/X _0809_/C VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0602__A2 _0597_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0888__A _0888_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_38 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_29_136 VSS VDD sky130_fd_sc_hd__fill_2
X_0739_ _0965_/A _0739_/B _0738_/X _0740_/C VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1024__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_172 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0841__A2 _0907_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0798__A _0924_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0964__C _0963_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_82 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_60 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_370 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0980__B _0930_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_301 VSS VDD sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X _1022_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XPHY_381 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0573_/A _0524_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1019__D _0558_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_18 VSS VDD sky130_fd_sc_hd__decap_4
X_1007_ _0809_/A _1007_/B _1007_/C _1008_/C VSS VDD sky130_fd_sc_hd__and3_4
XPHY_18 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_29 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_39 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_17 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0890__B _0901_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0823__A2 _0614_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_216 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1000__A2 _0749_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0784__C _0783_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_84 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0578__A1 _0512_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0750__A1 PAR_IN8[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0975__B _0971_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0991__A PAR_IN5[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0805__A2 _0730_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_194 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0569__A1 _0559_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_49 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_186 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_278 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_201 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_50 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_71 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_61 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_164 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0971__A1 PAR_IN7[28] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0986__A _0933_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_87 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_259 VSS VDD sky130_fd_sc_hd__fill_2
X_0987_ _0810_/A _0976_/X _0986_/X _0987_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0962__A1 PAR_IN7[8] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0896__A PAR_IN7[14] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0714__A1 PAR_IN3[27] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_259 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_278 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_189 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_82 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_267 VSS VDD sky130_fd_sc_hd__fill_1
X_0910_ _0976_/A _0901_/X _0910_/C _0910_/X VSS VDD sky130_fd_sc_hd__and3_4
X_0841_ PAR_IN8[10] _0907_/B _0615_/A _0844_/C VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0641__B1 _0640_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0772_ _0766_/X _0768_/X _0772_/C _0771_/X _0773_/C VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_45_3 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1027__D _0555_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_248 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_259 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0871__B1 _0870_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_229 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_95 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0926__A1 PAR_IN3[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_163 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0983__B _0994_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_218 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_207 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_0_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_281 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0917__A1 PAR_IN2[6] VSS VDD sky130_fd_sc_hd__diode_2
X_0755_ PAR_IN3[21] _0725_/X _0754_/X _0761_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_0824_ PAR_IN5[17] _0610_/B _0824_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_29_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_29 VSS VDD sky130_fd_sc_hd__fill_2
X_0686_ PAR_IN1[3] _0593_/B _0697_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0877__C _0877_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_17 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0893__B _0608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0853__B1 _0852_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_262 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0908__A1 PAR_IN2[22] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_159 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_83 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_211 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_295 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0978__B _0946_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0540_ _0530_/X _0534_/X _0540_/C _0540_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0697__C _0697_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_118 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0994__A PAR_IN6[4] VSS VDD sky130_fd_sc_hd__diode_2
X_1023_ _1023_/D COUNT[4] RESET _1020_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_0807_ PAR_IN7[25] _0689_/X _0806_/X _0807_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0738_ _0512_/X _0723_/X _0737_/X _0738_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__0888__B _0888_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0669_ _0619_/A _0946_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_52_162 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_129 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_118 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_302 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0826__B1 _0616_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1003__B1 _0616_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_247 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_269 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_382 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_82 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_195 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0989__A PAR_IN2[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_98 VSS VDD sky130_fd_sc_hd__fill_2
X_0523_ _0522_/X _0573_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_34_162 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_140 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_129 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_181 VSS VDD sky130_fd_sc_hd__fill_2
X_1006_ _1000_/X _1002_/X _1003_/X _1006_/D _1007_/C VSS VDD sky130_fd_sc_hd__or4_4
XPHY_19 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0899__A _0510_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_154 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0578__A2 _0577_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_232 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_221 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0975__C _0975_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0750__A2 _0677_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_287 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0991__B _0930_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_151 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0569__A2 _0567_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_190 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0512__A _0933_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_243 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_28 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_110 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_305 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_22_198 VSS VDD sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X _1020_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_45_235 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_83 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_169 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_110 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_176 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0971__A2 _0645_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_11 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0986__B _0986_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_268 VSS VDD sky130_fd_sc_hd__fill_2
X_0986_ _0933_/A _0986_/B _0985_/X _0986_/X VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_8_180 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0962__A2 _0689_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_17 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0896__B _0896_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0714__A2 _0635_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_257 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_293 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_290 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_238 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_216 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_205 VSS VDD sky130_fd_sc_hd__decap_4
X_0771_ PAR_IN7[29] _0706_/X _0770_/X _0771_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0840_ PAR_IN7[10] _0623_/A _0839_/X _0840_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0641__A1 PAR_IN8[31] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0997__A _0933_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_227 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_24_205 VSS VDD sky130_fd_sc_hd__decap_8
X_0969_ PAR_IN3[28] _0634_/X _0968_/X _0969_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_3_109 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1018__RESET_B RESET VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0871__A1 PAR_IN6[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_85 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_52 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0926__A2 _0634_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0610__A PAR_IN5[15] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_82 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_54 VSS VDD sky130_fd_sc_hd__fill_2
X_0685_ _1009_/A _0652_/Y _0684_/Y _0685_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0917__A2 _0699_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0823_ PAR_IN3[17] _0614_/X _0822_/X _0823_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_0754_ PAR_IN2[21] _0671_/B _0754_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0520__A _0810_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0877__D _0876_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0853__A1 PAR_IN2[26] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0908__A2 _0956_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1020__CLK _1020_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_149 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_138 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_300 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_52 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0605__A _0907_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_234 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_278 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0994__B _0994_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_105 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0532__B1 READY VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_182 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_138 VSS VDD sky130_fd_sc_hd__fill_2
X_1022_ _1022_/D COUNT[3] RESET _1022_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__0515__A COUNT[2] VSS VDD sky130_fd_sc_hd__diode_2
X_0806_ PAR_IN6[25] _0994_/B _0806_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0771__B1 _0770_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0668_ PAR_IN1[23] _0631_/X _0668_/X VSS VDD sky130_fd_sc_hd__or2_4
X_0737_ _0737_/A _0729_/X _0734_/X _0736_/X _0737_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0888__C _0888_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0599_ _0599_/A _0787_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_37_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_314 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_193 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0826__A1 PAR_IN4[17] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1003__A1 PAR_IN6[20] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_215 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_72 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_182 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_383 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_94 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0989__B _0946_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0522_ _0512_/X _0520_/X _0521_/Y _0522_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_20_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_174 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_160 VSS VDD sky130_fd_sc_hd__decap_12
X_1005_ PAR_IN4[20] _0692_/X _1004_/X _1006_/D VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__0899__B _0899_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0992__B1 _0991_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_177 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_144 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_111 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_200 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0975__D _0974_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_240 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0974__B1 _0973_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_180 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

