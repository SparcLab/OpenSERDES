/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */
/* With case-insensitive names (SPICE-compatible) */

module CLK_RECOVERY(
    inout vpwr,
    inout vgnd,
    input BB_IN,
    input CLK_IN,
    output CLK_OUT,
    output DATA_OUT,
    input RESET_N,
    input VDD,
    input VSS,
    input [21:0] SCAN_IN
);

wire _0719_ ;
wire _0892_ ;
wire _0472_ ;
wire _0052_ ;
wire _0528_ ;
wire _0108_ ;
wire _0281_ ;
wire _0757_ ;
wire _0337_ ;
wire _0090_ ;
wire _0566_ ;
wire _0146_ ;
wire _0795_ ;
wire _0375_ ;
wire _0184_ ;
wire _0889_ ;
wire _0469_ ;
wire _0049_ ;
wire _0698_ ;
wire _0278_ ;
wire _0910_ ;
wire _0087_ ;
wire clknet_1_0__leaf_clk_0_16 ;
wire _0813_ ;
wire _0622_ ;
wire _0202_ ;
wire _0851_ ;
wire _0431_ ;
wire _0011_ ;
wire _0907_ ;
wire _0660_ ;
wire _0240_ ;
wire _0716_ ;
wire _0525_ ;
wire _0105_ ;
wire _0754_ ;
wire _0334_ ;
wire _0563_ ;
wire _0143_ ;
wire _0619_ ;
wire _0792_ ;
wire _0372_ ;
wire _0848_ ;
wire _0428_ ;
wire _0008_ ;
wire BB_IN ;
wire _0181_ ;
wire _0657_ ;
wire _0237_ ;
wire _0886_ ;
wire _0466_ ;
wire _0046_ ;
wire _0695_ ;
wire _0275_ ;
wire _0084_ ;
wire \COUNT_BB_ONE[8]  ;
wire _0789_ ;
wire _0369_ ;
wire \COUNT_MIN[1]  ;
wire _0598_ ;
wire _0178_ ;
wire _0810_ ;
wire clknet_1_1__leaf_clk_0_32 ;
wire \COUNT_BB_ONE_MIN[4]  ;
wire _0904_ ;
wire _0713_ ;
wire _0522_ ;
wire _0102_ ;
wire _0751_ ;
wire _0331_ ;
wire _0807_ ;
wire _0560_ ;
wire _0140_ ;
wire _0616_ ;
wire _0845_ ;
wire _0425_ ;
wire _0005_ ;
wire _0654_ ;
wire _0234_ ;
wire \COUNT_BB_ZERO_MIN[0]  ;
wire \COUNT_BB_ZERO[5]  ;
wire _0883_ ;
wire _0463_ ;
wire _0043_ ;
wire _0519_ ;
wire _0692_ ;
wire _0272_ ;
wire _0748_ ;
wire _0328_ ;
wire _0081_ ;
wire _0557_ ;
wire _0137_ ;
wire _0786_ ;
wire _0366_ ;
wire _0595_ ;
wire _0175_ ;
wire _0689_ ;
wire _0269_ ;
wire _0901_ ;
wire _0498_ ;
wire _0078_ ;
wire _0710_ ;
wire clk_0_48 ;
wire _0804_ ;
wire _0613_ ;
wire \COUNT_BB_ZERO_MIN[10]  ;
wire _0842_ ;
wire _0422_ ;
wire _0002_ ;
wire \COUNT_MIN[8]  ;
wire _0651_ ;
wire _0231_ ;
wire _0707_ ;
wire _0880_ ;
wire _0460_ ;
wire _0040_ ;
wire _0516_ ;
wire _0745_ ;
wire _0325_ ;
wire _0554_ ;
wire _0134_ ;
wire _0783_ ;
wire _0363_ ;
wire _0839_ ;
wire _0419_ ;
wire _0592_ ;
wire _0172_ ;
wire _0648_ ;
wire _0228_ ;
wire _0877_ ;
wire _0457_ ;
wire _0037_ ;
wire \DIVISOR_COUNT[5]  ;
wire _0686_ ;
wire _0266_ ;
wire _0495_ ;
wire _0075_ ;
wire clk_0_16 ;
wire \COUNT_BB_ZERO_MIN[7]  ;
wire _0589_ ;
wire _0169_ ;
wire _0801_ ;
wire _0398_ ;
wire _0610_ ;
wire _0704_ ;
wire _0513_ ;
wire _0742_ ;
wire _0322_ ;
wire _0551_ ;
wire _0131_ ;
wire _0607_ ;
wire _0780_ ;
wire _0360_ ;
wire _0836_ ;
wire _0416_ ;
wire _0645_ ;
wire _0225_ ;
wire _0874_ ;
wire _0454_ ;
wire _0034_ ;
wire \COUNT_BB_ONE[3]  ;
wire _0683_ ;
wire _0263_ ;
wire _0739_ ;
wire _0319_ ;
wire _0492_ ;
wire _0072_ ;
wire _0548_ ;
wire _0128_ ;
wire _0777_ ;
wire _0357_ ;
wire _0586_ ;
wire _0166_ ;
wire _0395_ ;
wire _0489_ ;
wire _0069_ ;
wire _0701_ ;
wire _0298_ ;
wire _0510_ ;
wire _0604_ ;
wire \COUNT_BB_ZERO[0]  ;
wire _0833_ ;
wire _0413_ ;
wire _0642_ ;
wire _0222_ ;
wire _0871_ ;
wire _0451_ ;
wire _0031_ ;
wire _0507_ ;
wire _0680_ ;
wire _0260_ ;
wire _0736_ ;
wire _0316_ ;
wire _0545_ ;
wire _0125_ ;
wire clknet_1_0_0_clk_1_0 ;
wire _0774_ ;
wire _0354_ ;
wire _0583_ ;
wire _0163_ ;
wire _0639_ ;
wire _0219_ ;
wire _0392_ ;
wire _0868_ ;
wire _0448_ ;
wire _0028_ ;
wire _0677_ ;
wire _0257_ ;
wire _0486_ ;
wire _0066_ ;
wire _0295_ ;
wire _0389_ ;
wire \COUNT_MIN[3]  ;
wire _0601_ ;
wire _0198_ ;
wire _0830_ ;
wire _0410_ ;
wire \COUNT_BB_ONE_MIN[6]  ;
wire _0924_ ;
wire _0504_ ;
wire _0733_ ;
wire _0313_ ;
wire _0542_ ;
wire _0122_ ;
wire _0771_ ;
wire _0351_ ;
wire _0827_ ;
wire _0407_ ;
wire _0580_ ;
wire _0160_ ;
wire \DIVISOR_COUNT[0]  ;
wire _0636_ ;
wire _0216_ ;
wire _0865_ ;
wire _0445_ ;
wire _0025_ ;
wire _0674_ ;
wire _0254_ ;
wire \COUNT_BB_ZERO_MIN[2]  ;
wire \COUNT_BB_ZERO[7]  ;
wire _0483_ ;
wire _0063_ ;
wire _0539_ ;
wire _0119_ ;
wire _0292_ ;
wire _0768_ ;
wire _0348_ ;
wire _0577_ ;
wire _0157_ ;
wire N_CLK ;
wire _0386_ ;
wire VSS ;
wire _0195_ ;
wire _0289_ ;
wire _0921_ ;
wire _0501_ ;
wire _0098_ ;
wire _0730_ ;
wire _0310_ ;
wire _0824_ ;
wire _0404_ ;
wire _0633_ ;
wire _0213_ ;
wire clknet_1_1_0_clk_0_48 ;
wire _0862_ ;
wire _0442_ ;
wire _0022_ ;
wire _0918_ ;
wire _0671_ ;
wire _0251_ ;
wire _0727_ ;
wire _0307_ ;
wire _0480_ ;
wire _0060_ ;
wire _0536_ ;
wire _0116_ ;
wire \COUNT_BB_ZERO[10]  ;
wire _0765_ ;
wire _0345_ ;
wire clknet_1_1_0_clk_1_0 ;
wire _0574_ ;
wire _0154_ ;
wire _0383_ ;
wire _0859_ ;
wire _0439_ ;
wire _0019_ ;
wire clknet_0_clk_0_0 ;
wire _0192_ ;
wire _0668_ ;
wire _0248_ ;
wire _0897_ ;
wire _0477_ ;
wire _0057_ ;
wire \DIVISOR_COUNT[7]  ;
wire _0286_ ;
wire DATA_OUT ;
wire _0095_ ;
wire \COUNT_BB_ZERO_MIN[9]  ;
wire _0189_ ;
wire _0821_ ;
wire _0401_ ;
wire _0630_ ;
wire _0210_ ;
wire _0915_ ;
wire _0724_ ;
wire _0304_ ;
wire _0533_ ;
wire _0113_ ;
wire _0762_ ;
wire _0342_ ;
wire _0818_ ;
wire _0571_ ;
wire _0151_ ;
wire _0627_ ;
wire _0207_ ;
wire _0380_ ;
wire _0856_ ;
wire _0436_ ;
wire _0016_ ;
wire _0665_ ;
wire _0245_ ;
wire _0894_ ;
wire _0474_ ;
wire _0054_ ;
wire \COUNT_BB_ONE[5]  ;
wire _0283_ ;
wire _0759_ ;
wire _0339_ ;
wire _0092_ ;
wire _0568_ ;
wire _0148_ ;
wire \COUNT_BB_ONE_MIN[1]  ;
wire _0797_ ;
wire _0377_ ;
wire _0186_ ;
wire RESET_LIFTED_N ;
wire RESET_LIFTED_P ;
wire _0912_ ;
wire _0089_ ;
wire _0721_ ;
wire _0301_ ;
wire clknet_1_0__leaf_clk_0_32 ;
wire _0530_ ;
wire _0110_ ;
wire _0815_ ;
wire _0624_ ;
wire _0204_ ;
wire \COUNT_BB_ZERO[2]  ;
wire _0853_ ;
wire _0433_ ;
wire _0013_ ;
wire _0909_ ;
wire _0662_ ;
wire _0242_ ;
wire _0718_ ;
wire _0891_ ;
wire _0471_ ;
wire _0051_ ;
wire _0527_ ;
wire _0107_ ;
wire _0280_ ;
wire _0756_ ;
wire _0336_ ;
wire _0565_ ;
wire _0145_ ;
wire _0794_ ;
wire _0374_ ;
wire _0183_ ;
wire _0659_ ;
wire _0239_ ;
wire _0888_ ;
wire _0468_ ;
wire _0048_ ;
wire _0697_ ;
wire _0277_ ;
wire _0086_ ;
wire MULTIBIT_ZERO ;
wire _0812_ ;
wire \COUNT_MIN[5]  ;
wire _0621_ ;
wire _0201_ ;
wire _0850_ ;
wire _0430_ ;
wire _0010_ ;
wire \COUNT_BB_ONE_MIN[8]  ;
wire _0906_ ;
wire _0715_ ;
wire _0524_ ;
wire _0104_ ;
wire _0753_ ;
wire _0333_ ;
wire \COUNT_BB_ONE_MIN[10]  ;
wire _0809_ ;
wire _0562_ ;
wire _0142_ ;
wire _0618_ ;
wire _0791_ ;
wire _0371_ ;
wire _0847_ ;
wire _0427_ ;
wire _0007_ ;
wire _0180_ ;
wire \DIVISOR_COUNT[2]  ;
wire _0656_ ;
wire _0236_ ;
wire _0885_ ;
wire _0465_ ;
wire _0045_ ;
wire clknet_0_clk_0_48 ;
wire _0694_ ;
wire _0274_ ;
wire clk_0_0 ;
wire \COUNT_BB_ZERO_MIN[4]  ;
wire \COUNT_BB_ZERO[9]  ;
wire _0083_ ;
wire _0559_ ;
wire _0139_ ;
wire _0788_ ;
wire _0368_ ;
wire _0597_ ;
wire _0177_ ;
wire VDD ;
wire _0903_ ;
wire _0712_ ;
wire _0521_ ;
wire _0101_ ;
wire _0750_ ;
wire _0330_ ;
wire _0806_ ;
wire _0615_ ;
wire _0844_ ;
wire _0424_ ;
wire _0004_ ;
wire RESET_LIFTED ;
wire \COUNT_BB_ONE[0]  ;
wire _0653_ ;
wire _0233_ ;
wire _0709_ ;
wire _0882_ ;
wire _0462_ ;
wire _0042_ ;
wire clknet_0_clk_0_16 ;
wire _0518_ ;
wire _0691_ ;
wire _0271_ ;
wire _0747_ ;
wire _0327_ ;
wire _0080_ ;
wire _0556_ ;
wire _0136_ ;
wire _0785_ ;
wire _0365_ ;
wire _0594_ ;
wire _0174_ ;
wire _0879_ ;
wire _0459_ ;
wire _0039_ ;
wire _0688_ ;
wire _0268_ ;
wire _0900_ ;
wire _0497_ ;
wire _0077_ ;
wire \DIVISOR_COUNT[9]  ;
wire clk_0_32 ;
wire _0803_ ;
wire _0612_ ;
wire _0841_ ;
wire _0421_ ;
wire _0001_ ;
wire _0650_ ;
wire _0230_ ;
wire _0706_ ;
wire _0515_ ;
wire _0744_ ;
wire _0324_ ;
wire _0553_ ;
wire _0133_ ;
wire _0609_ ;
wire _0782_ ;
wire _0362_ ;
wire _0838_ ;
wire _0418_ ;
wire _0591_ ;
wire _0171_ ;
wire _0647_ ;
wire _0227_ ;
wire _0876_ ;
wire _0456_ ;
wire _0036_ ;
wire _0685_ ;
wire _0265_ ;
wire _0494_ ;
wire _0074_ ;
wire \COUNT_BB_ONE[7]  ;
wire _0779_ ;
wire _0359_ ;
wire \COUNT_MIN[0]  ;
wire _0588_ ;
wire _0168_ ;
wire _0800_ ;
wire \COUNT_BB_ONE_MIN[3]  ;
wire _0397_ ;
wire _0703_ ;
wire _0512_ ;
wire _0741_ ;
wire _0321_ ;
wire _0550_ ;
wire _0130_ ;
wire _0606_ ;
wire _0835_ ;
wire _0415_ ;
wire _0644_ ;
wire _0224_ ;
wire \COUNT_BB_ZERO[4]  ;
wire _0873_ ;
wire _0453_ ;
wire _0033_ ;
wire _0509_ ;
wire _0682_ ;
wire _0262_ ;
wire _0738_ ;
wire _0318_ ;
wire _0491_ ;
wire _0071_ ;
wire _0547_ ;
wire _0127_ ;
wire _0776_ ;
wire _0356_ ;
wire CLK_IN ;
wire _0585_ ;
wire _0165_ ;
wire _0394_ ;
wire _0679_ ;
wire _0259_ ;
wire _0488_ ;
wire _0068_ ;
wire _0700_ ;
wire _0297_ ;
wire _0603_ ;
wire _0832_ ;
wire _0412_ ;
wire \COUNT_MIN[7]  ;
wire _0641_ ;
wire _0221_ ;
wire _0870_ ;
wire _0450_ ;
wire _0030_ ;
wire _0506_ ;
wire _0735_ ;
wire _0315_ ;
wire _0544_ ;
wire _0124_ ;
wire _0773_ ;
wire _0353_ ;
wire _0829_ ;
wire _0409_ ;
wire _0582_ ;
wire _0162_ ;
wire _0638_ ;
wire _0218_ ;
wire _0391_ ;
wire _0867_ ;
wire _0447_ ;
wire _0027_ ;
wire \DIVISOR_COUNT[4]  ;
wire _0676_ ;
wire _0256_ ;
wire _0485_ ;
wire _0065_ ;
wire _0294_ ;
wire \COUNT_BB_ZERO_MIN[6]  ;
wire _0579_ ;
wire _0159_ ;
wire _0388_ ;
wire _0600_ ;
wire _0197_ ;
wire _0923_ ;
wire _0503_ ;
wire _0732_ ;
wire _0312_ ;
wire _0541_ ;
wire _0121_ ;
wire _0770_ ;
wire _0350_ ;
wire _0826_ ;
wire _0406_ ;
wire _0635_ ;
wire _0215_ ;
wire _0864_ ;
wire _0444_ ;
wire _0024_ ;
wire \COUNT_BB_ONE[2]  ;
wire _0673_ ;
wire _0253_ ;
wire _0729_ ;
wire _0309_ ;
wire _0482_ ;
wire _0062_ ;
wire _0538_ ;
wire _0118_ ;
wire _0291_ ;
wire _0767_ ;
wire _0347_ ;
wire _0576_ ;
wire _0156_ ;
wire _0385_ ;
wire _0194_ ;
wire _0899_ ;
wire _0479_ ;
wire _0059_ ;
wire _0288_ ;
wire _0920_ ;
wire _0500_ ;
wire _0097_ ;
wire _0823_ ;
wire _0403_ ;
wire _0632_ ;
wire _0212_ ;
wire _0861_ ;
wire _0441_ ;
wire _0021_ ;
wire _0917_ ;
wire _0670_ ;
wire _0250_ ;
wire _0726_ ;
wire _0306_ ;
wire _0535_ ;
wire _0115_ ;
wire clknet_1_0_0_clk_0_0 ;
wire _0764_ ;
wire _0344_ ;
wire _0573_ ;
wire _0153_ ;
wire _0629_ ;
wire _0209_ ;
wire _0382_ ;
wire _0858_ ;
wire _0438_ ;
wire _0018_ ;
wire _0191_ ;
wire _0667_ ;
wire _0247_ ;
wire _0896_ ;
wire _0476_ ;
wire _0056_ ;
wire _0285_ ;
wire _0094_ ;
wire \COUNT_BB_ONE[9]  ;
wire _0799_ ;
wire _0379_ ;
wire \COUNT_MIN[2]  ;
wire _0188_ ;
wire _0820_ ;
wire _0400_ ;
wire \COUNT_BB_ONE_MIN[5]  ;
wire _0914_ ;
wire _0723_ ;
wire _0303_ ;
wire _0532_ ;
wire _0112_ ;
wire RESET_N ;
wire _0761_ ;
wire _0341_ ;
wire _0817_ ;
wire _0570_ ;
wire _0150_ ;
wire _0626_ ;
wire _0206_ ;
wire CLK_OUT ;
wire _0855_ ;
wire _0435_ ;
wire _0015_ ;
wire _0664_ ;
wire _0244_ ;
wire \COUNT_BB_ZERO_MIN[1]  ;
wire \COUNT_BB_ZERO[6]  ;
wire _0893_ ;
wire _0473_ ;
wire _0053_ ;
wire _0529_ ;
wire _0109_ ;
wire _0282_ ;
wire _0758_ ;
wire _0338_ ;
wire _0091_ ;
wire _0567_ ;
wire _0147_ ;
wire _0796_ ;
wire _0376_ ;
wire _0185_ ;
wire _0699_ ;
wire _0279_ ;
wire _0911_ ;
wire _0088_ ;
wire _0720_ ;
wire _0300_ ;
wire _0814_ ;
wire _0623_ ;
wire _0203_ ;
wire _0852_ ;
wire _0432_ ;
wire _0012_ ;
wire \COUNT_MIN[9]  ;
wire _0908_ ;
wire _0661_ ;
wire _0241_ ;
wire _0717_ ;
wire _0890_ ;
wire _0470_ ;
wire _0050_ ;
wire _0526_ ;
wire _0106_ ;
wire _0755_ ;
wire _0335_ ;
wire clknet_1_1_0_clk_0_0 ;
wire _0564_ ;
wire _0144_ ;
wire _0793_ ;
wire _0373_ ;
wire ZERO_CHECKED ;
wire _0849_ ;
wire _0429_ ;
wire _0009_ ;
wire _0182_ ;
wire _0658_ ;
wire _0238_ ;
wire _0887_ ;
wire _0467_ ;
wire _0047_ ;
wire \DIVISOR_COUNT[6]  ;
wire _0696_ ;
wire _0276_ ;
wire _0085_ ;
wire \COUNT_BB_ZERO_MIN[8]  ;
wire _0599_ ;
wire _0179_ ;
wire _0811_ ;
wire _0620_ ;
wire _0200_ ;
wire _0905_ ;
wire _0714_ ;
wire _0523_ ;
wire _0103_ ;
wire _0752_ ;
wire _0332_ ;
wire _0808_ ;
wire _0561_ ;
wire _0141_ ;
wire _0617_ ;
wire _0790_ ;
wire _0370_ ;
wire _0846_ ;
wire _0426_ ;
wire _0006_ ;
wire _0655_ ;
wire _0235_ ;
wire _0884_ ;
wire _0464_ ;
wire _0044_ ;
wire \COUNT_BB_ONE[4]  ;
wire clknet_0_clk_0_32 ;
wire _0693_ ;
wire _0273_ ;
wire _0749_ ;
wire _0329_ ;
wire _0082_ ;
wire _0558_ ;
wire _0138_ ;
wire \COUNT_BB_ONE_MIN[0]  ;
wire _0787_ ;
wire _0367_ ;
wire _0596_ ;
wire _0176_ ;
wire clknet_1_1__leaf_clk_0_16 ;
wire _0902_ ;
wire _0499_ ;
wire _0079_ ;
wire _0711_ ;
wire _0520_ ;
wire _0100_ ;
wire _0805_ ;
wire _0614_ ;
wire \COUNT_BB_ZERO[1]  ;
wire _0843_ ;
wire _0423_ ;
wire _0003_ ;
wire _0652_ ;
wire _0232_ ;
wire _0708_ ;
wire _0881_ ;
wire _0461_ ;
wire _0041_ ;
wire _0517_ ;
wire _0690_ ;
wire _0270_ ;
wire _0746_ ;
wire _0326_ ;
wire _0555_ ;
wire _0135_ ;
wire _0784_ ;
wire _0364_ ;
wire _0593_ ;
wire _0173_ ;
wire _0649_ ;
wire _0229_ ;
wire _0878_ ;
wire _0458_ ;
wire _0038_ ;
wire _0687_ ;
wire _0267_ ;
wire _0496_ ;
wire _0076_ ;
wire _0802_ ;
wire _0399_ ;
wire \COUNT_MIN[4]  ;
wire _0611_ ;
wire _0840_ ;
wire _0420_ ;
wire _0000_ ;
wire \COUNT_BB_ONE_MIN[7]  ;
wire _0705_ ;
wire _0514_ ;
wire _0743_ ;
wire _0323_ ;
wire _0552_ ;
wire _0132_ ;
wire MULTIBIT_ONE ;
wire _0608_ ;
wire _0781_ ;
wire _0361_ ;
wire _0837_ ;
wire _0417_ ;
wire _0590_ ;
wire _0170_ ;
wire \DIVISOR_COUNT[1]  ;
wire _0646_ ;
wire _0226_ ;
wire _0875_ ;
wire _0455_ ;
wire _0035_ ;
wire _0684_ ;
wire _0264_ ;
wire \COUNT_BB_ZERO_MIN[3]  ;
wire \COUNT_BB_ZERO[8]  ;
wire _0493_ ;
wire _0073_ ;
wire _0549_ ;
wire _0129_ ;
wire _0778_ ;
wire _0358_ ;
wire _0587_ ;
wire _0167_ ;
wire _0396_ ;
wire _0702_ ;
wire _0299_ ;
wire _0511_ ;
wire _0740_ ;
wire _0320_ ;
wire _0605_ ;
wire _0834_ ;
wire _0414_ ;
wire _0643_ ;
wire _0223_ ;
wire P_CLK ;
wire _0872_ ;
wire _0452_ ;
wire _0032_ ;
wire _0508_ ;
wire _0681_ ;
wire _0261_ ;
wire _0737_ ;
wire _0317_ ;
wire _0490_ ;
wire _0070_ ;
wire _0546_ ;
wire _0126_ ;
wire _0775_ ;
wire _0355_ ;
wire _0584_ ;
wire _0164_ ;
wire _0393_ ;
wire _0869_ ;
wire _0449_ ;
wire _0029_ ;
wire clknet_0_clk_1_0 ;
wire _0678_ ;
wire _0258_ ;
wire _0487_ ;
wire _0067_ ;
wire \DIVISOR_COUNT[8]  ;
wire _0296_ ;
wire _0602_ ;
wire _0199_ ;
wire _0831_ ;
wire _0411_ ;
wire _0640_ ;
wire _0220_ ;
wire _0505_ ;
wire _0734_ ;
wire _0314_ ;
wire _0543_ ;
wire _0123_ ;
wire _0772_ ;
wire _0352_ ;
wire _0828_ ;
wire _0408_ ;
wire _0581_ ;
wire _0161_ ;
wire _0637_ ;
wire _0217_ ;
wire _0390_ ;
wire _0866_ ;
wire _0446_ ;
wire _0026_ ;
wire _0675_ ;
wire _0255_ ;
wire _0484_ ;
wire _0064_ ;
wire \COUNT_BB_ONE[6]  ;
wire _0293_ ;
wire _0769_ ;
wire _0349_ ;
wire \DIVISOR_COUNT[10]  ;
wire _0578_ ;
wire _0158_ ;
wire \COUNT_BB_ONE_MIN[2]  ;
wire _0387_ ;
wire _0196_ ;
wire _0922_ ;
wire _0502_ ;
wire _0099_ ;
wire _0731_ ;
wire _0311_ ;
wire _0540_ ;
wire _0120_ ;
wire _0825_ ;
wire _0405_ ;
wire _0634_ ;
wire _0214_ ;
wire \COUNT_BB_ZERO[3]  ;
wire _0863_ ;
wire _0443_ ;
wire _0023_ ;
wire _0919_ ;
wire _0672_ ;
wire _0252_ ;
wire _0728_ ;
wire _0308_ ;
wire _0481_ ;
wire _0061_ ;
wire _0537_ ;
wire _0117_ ;
wire _0290_ ;
wire _0766_ ;
wire _0346_ ;
wire _0575_ ;
wire _0155_ ;
wire _0384_ ;
wire _0193_ ;
wire _0669_ ;
wire _0249_ ;
wire _0898_ ;
wire _0478_ ;
wire _0058_ ;
wire _0287_ ;
wire _0096_ ;
wire \COUNT_BB_ONE[10]  ;
wire _0822_ ;
wire _0402_ ;
wire \COUNT_MIN[6]  ;
wire _0631_ ;
wire _0211_ ;
wire _0860_ ;
wire _0440_ ;
wire _0020_ ;
wire \COUNT_BB_ONE_MIN[9]  ;
wire _0916_ ;
wire _0725_ ;
wire _0305_ ;
wire _0534_ ;
wire _0114_ ;
wire _0763_ ;
wire _0343_ ;
wire _0819_ ;
wire _0572_ ;
wire _0152_ ;
wire _0628_ ;
wire _0208_ ;
wire _0381_ ;
wire _0857_ ;
wire _0437_ ;
wire _0017_ ;
wire _0190_ ;
wire \DIVISOR_COUNT[3]  ;
wire _0666_ ;
wire _0246_ ;
wire _0895_ ;
wire _0475_ ;
wire _0055_ ;
wire _0284_ ;
wire clk_1_0 ;
wire \COUNT_BB_ZERO_MIN[5]  ;
wire _0093_ ;
wire _0569_ ;
wire _0149_ ;
wire _0798_ ;
wire _0378_ ;
wire ONE_CHECKED ;
wire clknet_1_0_0_clk_0_48 ;
wire _0187_ ;
wire _0913_ ;
wire _0722_ ;
wire _0302_ ;
wire _0531_ ;
wire _0111_ ;
wire _0760_ ;
wire _0340_ ;
wire _0816_ ;
wire [21:0] SCAN_IN ;
wire _0625_ ;
wire _0205_ ;
wire _0854_ ;
wire _0434_ ;
wire _0014_ ;
wire \COUNT_BB_ONE[1]  ;
wire _0663_ ;
wire _0243_ ;

sky130_fd_sc_hd__inv_8 _0925_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(ONE_CHECKED),
    .Y(_0144_)
);

sky130_fd_sc_hd__inv_8 _0926_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(P_CLK),
    .Y(_0145_)
);

sky130_fd_sc_hd__a2bb2o_4 _0927_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0144_),
    .A2_N(_0145_),
    .B1(ZERO_CHECKED),
    .B2(_0145_),
    .X(_0146_)
);

sky130_fd_sc_hd__inv_8 _0928_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[9] ),
    .Y(_0147_)
);

sky130_fd_sc_hd__or3_4 _0929_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[0] ),
    .B(\COUNT_MIN[1] ),
    .C(\COUNT_MIN[2] ),
    .X(_0148_)
);

sky130_fd_sc_hd__or2_4 _0930_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[3] ),
    .B(_0148_),
    .X(_0149_)
);

sky130_fd_sc_hd__or2_4 _0931_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[4] ),
    .B(_0149_),
    .X(_0150_)
);

sky130_fd_sc_hd__or2_4 _0932_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[5] ),
    .B(_0150_),
    .X(_0151_)
);

sky130_fd_sc_hd__or2_4 _0933_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[6] ),
    .B(_0151_),
    .X(_0152_)
);

sky130_fd_sc_hd__or2_4 _0934_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[7] ),
    .B(_0152_),
    .X(_0153_)
);

sky130_fd_sc_hd__or2_4 _0935_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[8] ),
    .B(_0153_),
    .X(_0154_)
);

sky130_fd_sc_hd__inv_8 _0936_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0154_),
    .Y(_0155_)
);

sky130_fd_sc_hd__or2_4 _0937_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[9] ),
    .B(_0154_),
    .X(_0156_)
);

sky130_fd_sc_hd__o21a_4 _0938_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0147_),
    .A2(_0155_),
    .B1(_0156_),
    .X(_0157_)
);

sky130_fd_sc_hd__and2_4 _0939_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[9] ),
    .B(_0157_),
    .X(_0158_)
);

sky130_fd_sc_hd__or2_4 _0940_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[9] ),
    .B(_0157_),
    .X(_0159_)
);

sky130_fd_sc_hd__buf_1 _0941_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0159_),
    .X(_0160_)
);

sky130_fd_sc_hd__inv_8 _0942_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .Y(_0161_)
);

sky130_fd_sc_hd__inv_8 _0943_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[4] ),
    .Y(_0162_)
);

sky130_fd_sc_hd__buf_1 _0944_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0162_),
    .X(_0163_)
);

sky130_fd_sc_hd__a21bo_4 _0945_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[4] ),
    .A2(_0149_),
    .B1_N(_0150_),
    .X(_0164_)
);

sky130_fd_sc_hd__inv_8 _0946_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[5] ),
    .Y(_0165_)
);

sky130_fd_sc_hd__a21bo_4 _0947_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[5] ),
    .A2(_0150_),
    .B1_N(_0151_),
    .X(_0166_)
);

sky130_fd_sc_hd__and2_4 _0948_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0165_),
    .B(_0166_),
    .X(_0167_)
);

sky130_fd_sc_hd__buf_1 _0949_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0167_),
    .X(_0168_)
);

sky130_fd_sc_hd__buf_1 _0950_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0165_),
    .X(_0169_)
);

sky130_fd_sc_hd__or2_4 _0951_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0162_),
    .B(_0164_),
    .X(_0170_)
);

sky130_fd_sc_hd__o21ai_4 _0952_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0169_),
    .A2(_0166_),
    .B1(_0170_),
    .Y(_0171_)
);

sky130_fd_sc_hd__a211o_4 _0953_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0163_),
    .A2(_0164_),
    .B1(_0168_),
    .C1(_0171_),
    .X(_0172_)
);

sky130_fd_sc_hd__a21boi_4 _0954_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[3] ),
    .A2(_0148_),
    .B1_N(_0149_),
    .Y(_0173_)
);

sky130_fd_sc_hd__or2_4 _0955_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[3] ),
    .B(_0173_),
    .X(_0174_)
);

sky130_fd_sc_hd__buf_1 _0956_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0174_),
    .X(_0175_)
);

sky130_fd_sc_hd__inv_8 _0957_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0175_),
    .Y(_0176_)
);

sky130_fd_sc_hd__inv_8 _0958_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[2] ),
    .Y(_0177_)
);

sky130_fd_sc_hd__inv_8 _0959_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[0] ),
    .Y(_0178_)
);

sky130_fd_sc_hd__inv_8 _0960_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[1] ),
    .Y(_0179_)
);

sky130_fd_sc_hd__and2_4 _0961_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0178_),
    .B(_0179_),
    .X(_0180_)
);

sky130_fd_sc_hd__o21a_4 _0962_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0177_),
    .A2(_0180_),
    .B1(_0148_),
    .X(_0181_)
);

sky130_fd_sc_hd__nor2_4 _0963_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[2] ),
    .B(_0181_),
    .Y(_0182_)
);

sky130_fd_sc_hd__inv_8 _0964_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[0] ),
    .Y(_0183_)
);

sky130_fd_sc_hd__inv_8 _0965_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[1] ),
    .Y(_0184_)
);

sky130_fd_sc_hd__a21o_4 _0966_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[0] ),
    .A2(\COUNT_MIN[1] ),
    .B1(_0180_),
    .X(_0185_)
);

sky130_fd_sc_hd__nor2_4 _0967_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0184_),
    .B(_0185_),
    .Y(_0186_)
);

sky130_fd_sc_hd__and2_4 _0968_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0184_),
    .B(_0185_),
    .X(_0187_)
);

sky130_fd_sc_hd__a211o_4 _0969_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0183_),
    .A2(_0178_),
    .B1(_0186_),
    .C1(_0187_),
    .X(_0188_)
);

sky130_fd_sc_hd__a211o_4 _0970_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\DIVISOR_COUNT[0] ),
    .A2(\COUNT_MIN[0] ),
    .B1(_0182_),
    .C1(_0188_),
    .X(_0189_)
);

sky130_fd_sc_hd__a22oi_4 _0971_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\DIVISOR_COUNT[3] ),
    .A2(_0173_),
    .B1(\DIVISOR_COUNT[2] ),
    .B2(_0181_),
    .Y(_0190_)
);

sky130_fd_sc_hd__inv_8 _0972_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0190_),
    .Y(_0191_)
);

sky130_fd_sc_hd__inv_8 _0973_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[7] ),
    .Y(_0192_)
);

sky130_fd_sc_hd__buf_1 _0974_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0192_),
    .X(_0193_)
);

sky130_fd_sc_hd__a21bo_4 _0975_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[7] ),
    .A2(_0152_),
    .B1_N(_0153_),
    .X(_0194_)
);

sky130_fd_sc_hd__nor2_4 _0976_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0193_),
    .B(_0194_),
    .Y(_0195_)
);

sky130_fd_sc_hd__or4_4 _0977_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0176_),
    .B(_0189_),
    .C(_0191_),
    .D(_0195_),
    .X(_0196_)
);

sky130_fd_sc_hd__inv_8 _0978_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[6] ),
    .Y(_0197_)
);

sky130_fd_sc_hd__a21bo_4 _0979_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[6] ),
    .A2(_0151_),
    .B1_N(_0152_),
    .X(_0198_)
);

sky130_fd_sc_hd__nor2_4 _0980_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0197_),
    .B(_0198_),
    .Y(_0199_)
);

sky130_fd_sc_hd__and2_4 _0981_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0192_),
    .B(_0194_),
    .X(_0200_)
);

sky130_fd_sc_hd__a211o_4 _0982_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0197_),
    .A2(_0198_),
    .B1(_0199_),
    .C1(_0200_),
    .X(_0201_)
);

sky130_fd_sc_hd__or2_4 _0983_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[10] ),
    .B(_0156_),
    .X(_0202_)
);

sky130_fd_sc_hd__buf_1 _0984_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0202_),
    .X(_0203_)
);

sky130_fd_sc_hd__inv_8 _0985_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0203_),
    .Y(_0204_)
);

sky130_fd_sc_hd__or4_4 _0986_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0172_),
    .B(_0196_),
    .C(_0201_),
    .D(_0204_),
    .X(_0205_)
);

sky130_fd_sc_hd__buf_1 _0987_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[10] ),
    .X(_0206_)
);

sky130_fd_sc_hd__inv_8 _0988_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[8] ),
    .Y(_0207_)
);

sky130_fd_sc_hd__buf_1 _0989_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0207_),
    .X(_0208_)
);

sky130_fd_sc_hd__a21o_4 _0990_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[8] ),
    .A2(_0153_),
    .B1(_0155_),
    .X(_0209_)
);

sky130_fd_sc_hd__nor2_4 _0991_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0208_),
    .B(_0209_),
    .Y(_0210_)
);

sky130_fd_sc_hd__and2_4 _0992_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0207_),
    .B(_0209_),
    .X(_0211_)
);

sky130_fd_sc_hd__buf_1 _0993_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0211_),
    .X(_0212_)
);

sky130_fd_sc_hd__a211o_4 _0994_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0206_),
    .A2(_0156_),
    .B1(_0210_),
    .C1(_0212_),
    .X(_0213_)
);

sky130_fd_sc_hd__nor4_4 _0995_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0158_),
    .B(_0161_),
    .C(_0205_),
    .D(_0213_),
    .Y(_0214_)
);

sky130_fd_sc_hd__or2_4 _0996_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0146_),
    .B(_0214_),
    .X(_0215_)
);

sky130_fd_sc_hd__buf_1 _0997_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0215_),
    .X(_0216_)
);

sky130_fd_sc_hd__inv_8 _0998_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0216_),
    .Y(_0217_)
);

sky130_fd_sc_hd__buf_1 _0999_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0183_),
    .X(_0218_)
);

sky130_fd_sc_hd__inv_8 _1000_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0212_),
    .Y(_0219_)
);

sky130_fd_sc_hd__inv_8 _1001_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0201_),
    .Y(_0220_)
);

sky130_fd_sc_hd__o21a_4 _1002_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0184_),
    .A2(_0185_),
    .B1(_0188_),
    .X(_0221_)
);

sky130_fd_sc_hd__o21ai_4 _1003_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0182_),
    .A2(_0221_),
    .B1(_0190_),
    .Y(_0222_)
);

sky130_fd_sc_hd__inv_8 _1004_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0172_),
    .Y(_0223_)
);

sky130_fd_sc_hd__inv_8 _1005_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0168_),
    .Y(_0224_)
);

sky130_fd_sc_hd__a32o_4 _1006_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0175_),
    .A2(_0222_),
    .A3(_0223_),
    .B1(_0224_),
    .B2(_0171_),
    .X(_0225_)
);

sky130_fd_sc_hd__nor3_4 _1007_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0197_),
    .B(_0198_),
    .C(_0200_),
    .Y(_0226_)
);

sky130_fd_sc_hd__a211o_4 _1008_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0220_),
    .A2(_0225_),
    .B1(_0195_),
    .C1(_0226_),
    .X(_0227_)
);

sky130_fd_sc_hd__a211o_4 _1009_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0219_),
    .A2(_0227_),
    .B1(_0210_),
    .C1(_0158_),
    .X(_0228_)
);

sky130_fd_sc_hd__a32o_4 _1010_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0203_),
    .A2(_0160_),
    .A3(_0228_),
    .B1(_0206_),
    .B2(_0156_),
    .X(_0229_)
);

sky130_fd_sc_hd__or2_4 _1011_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0218_),
    .B(_0229_),
    .X(_0230_)
);

sky130_fd_sc_hd__inv_8 _1012_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0229_),
    .Y(_0231_)
);

sky130_fd_sc_hd__or2_4 _1013_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[0] ),
    .B(_0231_),
    .X(_0232_)
);

sky130_fd_sc_hd__and3_4 _1014_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0217_),
    .B(_0230_),
    .C(_0232_),
    .X(_0055_)
);

sky130_fd_sc_hd__buf_1 _1015_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0184_),
    .X(_0233_)
);

sky130_fd_sc_hd__or3_4 _1016_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0218_),
    .B(_0233_),
    .C(_0229_),
    .X(_0234_)
);

sky130_fd_sc_hd__nand2_4 _1017_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0233_),
    .B(_0230_),
    .Y(_0235_)
);

sky130_fd_sc_hd__and3_4 _1018_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0217_),
    .B(_0234_),
    .C(_0235_),
    .X(_0057_)
);

sky130_fd_sc_hd__inv_8 _1019_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[2] ),
    .Y(_0236_)
);

sky130_fd_sc_hd__or4_4 _1020_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0218_),
    .B(_0233_),
    .C(_0236_),
    .D(_0229_),
    .X(_0237_)
);

sky130_fd_sc_hd__nand2_4 _1021_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0236_),
    .B(_0234_),
    .Y(_0238_)
);

sky130_fd_sc_hd__and3_4 _1022_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0217_),
    .B(_0237_),
    .C(_0238_),
    .X(_0058_)
);

sky130_fd_sc_hd__inv_8 _1023_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[3] ),
    .Y(_0239_)
);

sky130_fd_sc_hd__nand2_4 _1024_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0239_),
    .B(_0237_),
    .Y(_0240_)
);

sky130_fd_sc_hd__or2_4 _1025_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0239_),
    .B(_0237_),
    .X(_0241_)
);

sky130_fd_sc_hd__and3_4 _1026_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0217_),
    .B(_0240_),
    .C(_0241_),
    .X(_0059_)
);

sky130_fd_sc_hd__or2_4 _1027_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0239_),
    .B(_0163_),
    .X(_0242_)
);

sky130_fd_sc_hd__or4_4 _1028_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0218_),
    .B(_0184_),
    .C(_0236_),
    .D(_0242_),
    .X(_0243_)
);

sky130_fd_sc_hd__inv_8 _1029_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0243_),
    .Y(_0244_)
);

sky130_fd_sc_hd__a21o_4 _1030_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0231_),
    .A2(_0244_),
    .B1(_0216_),
    .X(_0245_)
);

sky130_fd_sc_hd__a21oi_4 _1031_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0163_),
    .A2(_0241_),
    .B1(_0245_),
    .Y(_0060_)
);

sky130_fd_sc_hd__buf_1 _1032_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0216_),
    .X(_0246_)
);

sky130_fd_sc_hd__or2_4 _1033_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[5] ),
    .B(_0244_),
    .X(_0247_)
);

sky130_fd_sc_hd__or2_4 _1034_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0169_),
    .B(_0243_),
    .X(_0248_)
);

sky130_fd_sc_hd__buf_1 _1035_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0229_),
    .X(_0249_)
);

sky130_fd_sc_hd__a21oi_4 _1036_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0247_),
    .A2(_0248_),
    .B1(_0249_),
    .Y(_0250_)
);

sky130_fd_sc_hd__nor2_4 _1037_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0231_),
    .B(_0214_),
    .Y(_0251_)
);

sky130_fd_sc_hd__and2_4 _1038_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0169_),
    .B(_0251_),
    .X(_0252_)
);

sky130_fd_sc_hd__nor3_4 _1039_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0246_),
    .B(_0250_),
    .C(_0252_),
    .Y(_0061_)
);

sky130_fd_sc_hd__buf_1 _1040_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0197_),
    .X(_0253_)
);

sky130_fd_sc_hd__or2_4 _1041_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0249_),
    .B(_0248_),
    .X(_0254_)
);

sky130_fd_sc_hd__a21oi_4 _1042_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0253_),
    .A2(_0254_),
    .B1(_0246_),
    .Y(_0255_)
);

sky130_fd_sc_hd__o21a_4 _1043_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0253_),
    .A2(_0254_),
    .B1(_0255_),
    .X(_0062_)
);

sky130_fd_sc_hd__or2_4 _1044_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0253_),
    .B(_0248_),
    .X(_0256_)
);

sky130_fd_sc_hd__or2_4 _1045_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0193_),
    .B(_0256_),
    .X(_0257_)
);

sky130_fd_sc_hd__a21boi_4 _1046_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0193_),
    .A2(_0256_),
    .B1_N(_0257_),
    .Y(_0258_)
);

sky130_fd_sc_hd__nor2_4 _1047_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0249_),
    .B(_0258_),
    .Y(_0259_)
);

sky130_fd_sc_hd__and2_4 _1048_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0193_),
    .B(_0251_),
    .X(_0260_)
);

sky130_fd_sc_hd__nor3_4 _1049_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0246_),
    .B(_0259_),
    .C(_0260_),
    .Y(_0063_)
);

sky130_fd_sc_hd__or2_4 _1050_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0249_),
    .B(_0257_),
    .X(_0261_)
);

sky130_fd_sc_hd__a21oi_4 _1051_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0208_),
    .A2(_0261_),
    .B1(_0246_),
    .Y(_0262_)
);

sky130_fd_sc_hd__o21a_4 _1052_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0208_),
    .A2(_0261_),
    .B1(_0262_),
    .X(_0064_)
);

sky130_fd_sc_hd__inv_8 _1053_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\DIVISOR_COUNT[9] ),
    .Y(_0263_)
);

sky130_fd_sc_hd__or2_4 _1054_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0208_),
    .B(_0257_),
    .X(_0264_)
);

sky130_fd_sc_hd__buf_1 _1055_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0264_),
    .X(_0265_)
);

sky130_fd_sc_hd__xor2_4 _1056_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0263_),
    .B(_0265_),
    .X(_0266_)
);

sky130_fd_sc_hd__nor2_4 _1057_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0249_),
    .B(_0266_),
    .Y(_0267_)
);

sky130_fd_sc_hd__and2_4 _1058_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0263_),
    .B(_0251_),
    .X(_0268_)
);

sky130_fd_sc_hd__nor3_4 _1059_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0246_),
    .B(_0267_),
    .C(_0268_),
    .Y(_0065_)
);

sky130_fd_sc_hd__nor3_4 _1060_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0263_),
    .B(_0265_),
    .C(_0251_),
    .Y(_0269_)
);

sky130_fd_sc_hd__nor2_4 _1061_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0206_),
    .B(_0269_),
    .Y(_0270_)
);

sky130_fd_sc_hd__and2_4 _1062_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0206_),
    .B(_0269_),
    .X(_0271_)
);

sky130_fd_sc_hd__nor3_4 _1063_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0146_),
    .B(_0270_),
    .C(_0271_),
    .Y(_0056_)
);

sky130_fd_sc_hd__buf_1 _1064_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(P_CLK),
    .X(_0272_)
);

sky130_fd_sc_hd__inv_8 _1065_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(ZERO_CHECKED),
    .Y(_0273_)
);

sky130_fd_sc_hd__nor2_4 _1066_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0273_),
    .B(CLK_OUT),
    .Y(_0274_)
);

sky130_fd_sc_hd__and2_4 _1067_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0239_),
    .B(\COUNT_MIN[4] ),
    .X(_0275_)
);

sky130_fd_sc_hd__and2_4 _1068_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[5] ),
    .B(_0163_),
    .X(_0276_)
);

sky130_fd_sc_hd__a211o_4 _1069_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[7] ),
    .A2(_0253_),
    .B1(_0275_),
    .C1(_0276_),
    .X(_0277_)
);

sky130_fd_sc_hd__or2_4 _1070_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[5] ),
    .B(_0163_),
    .X(_0278_)
);

sky130_fd_sc_hd__o21ai_4 _1071_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[6] ),
    .A2(_0169_),
    .B1(_0278_),
    .Y(_0279_)
);

sky130_fd_sc_hd__a2bb2o_4 _1072_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(\COUNT_MIN[7] ),
    .A2_N(_0253_),
    .B1(_0193_),
    .B2(\COUNT_MIN[8] ),
    .X(_0280_)
);

sky130_fd_sc_hd__a2bb2o_4 _1073_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(\COUNT_MIN[3] ),
    .A2_N(_0236_),
    .B1(\COUNT_MIN[3] ),
    .B2(_0236_),
    .X(_0281_)
);

sky130_fd_sc_hd__a2bb2o_4 _1074_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0233_),
    .A2_N(\COUNT_MIN[2] ),
    .B1(\COUNT_MIN[6] ),
    .B2(_0169_),
    .X(_0282_)
);

sky130_fd_sc_hd__or4_4 _1075_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0279_),
    .B(_0280_),
    .C(_0281_),
    .D(_0282_),
    .X(_0283_)
);

sky130_fd_sc_hd__inv_8 _1076_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_MIN[8] ),
    .Y(_0284_)
);

sky130_fd_sc_hd__a211o_4 _1077_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\DIVISOR_COUNT[7] ),
    .A2(_0284_),
    .B1(\DIVISOR_COUNT[9] ),
    .C1(_0206_),
    .X(_0285_)
);

sky130_fd_sc_hd__a2bb2o_4 _1078_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0239_),
    .A2_N(\COUNT_MIN[4] ),
    .B1(_0233_),
    .B2(\COUNT_MIN[2] ),
    .X(_0286_)
);

sky130_fd_sc_hd__o22a_4 _1079_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_MIN[9] ),
    .A2(\DIVISOR_COUNT[8] ),
    .B1(_0147_),
    .B2(_0208_),
    .X(_0287_)
);

sky130_fd_sc_hd__o22a_4 _1080_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\DIVISOR_COUNT[0] ),
    .A2(\COUNT_MIN[1] ),
    .B1(_0218_),
    .B2(_0179_),
    .X(_0288_)
);

sky130_fd_sc_hd__or4_4 _1081_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0285_),
    .B(_0286_),
    .C(_0287_),
    .D(_0288_),
    .X(_0289_)
);

sky130_fd_sc_hd__nor4_4 _1082_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0277_),
    .B(_0283_),
    .C(_0289_),
    .D(_0214_),
    .Y(_0290_)
);

sky130_fd_sc_hd__xnor2_4 _1083_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(CLK_OUT),
    .B(_0290_),
    .Y(_0291_)
);

sky130_fd_sc_hd__and2_4 _1084_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0273_),
    .B(_0291_),
    .X(_0292_)
);

sky130_fd_sc_hd__and2_4 _1085_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0144_),
    .B(_0291_),
    .X(_0293_)
);

sky130_fd_sc_hd__buf_1 _1086_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(P_CLK),
    .X(_0294_)
);

sky130_fd_sc_hd__o21ai_4 _1087_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0144_),
    .A2(CLK_OUT),
    .B1(_0294_),
    .Y(_0295_)
);

sky130_fd_sc_hd__o32ai_4 _1088_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0272_),
    .A2(_0274_),
    .A3(_0292_),
    .B1(_0293_),
    .B2(_0295_),
    .Y(_0000_)
);

sky130_fd_sc_hd__buf_1 _1089_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[1] ),
    .X(_0296_)
);

sky130_fd_sc_hd__or2_4 _1090_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0296_),
    .B(\COUNT_BB_ONE_MIN[0] ),
    .X(_0297_)
);

sky130_fd_sc_hd__inv_8 _1091_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[1] ),
    .Y(_0298_)
);

sky130_fd_sc_hd__inv_8 _1092_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[0] ),
    .Y(_0299_)
);

sky130_fd_sc_hd__or2_4 _1093_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0298_),
    .B(_0299_),
    .X(_0300_)
);

sky130_fd_sc_hd__buf_1 _1094_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[1] ),
    .X(_0301_)
);

sky130_fd_sc_hd__or2_4 _1095_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0301_),
    .B(\COUNT_BB_ZERO_MIN[0] ),
    .X(_0302_)
);

sky130_fd_sc_hd__inv_8 _1096_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[1] ),
    .Y(_0303_)
);

sky130_fd_sc_hd__buf_1 _1097_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0303_),
    .X(_0304_)
);

sky130_fd_sc_hd__inv_8 _1098_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[0] ),
    .Y(_0305_)
);

sky130_fd_sc_hd__buf_1 _1099_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0305_),
    .X(_0306_)
);

sky130_fd_sc_hd__buf_1 _1100_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0145_),
    .X(_0307_)
);

sky130_fd_sc_hd__o21a_4 _1101_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0304_),
    .A2(_0306_),
    .B1(_0307_),
    .X(_0308_)
);

sky130_fd_sc_hd__a32oi_4 _1102_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0272_),
    .A2(_0297_),
    .A3(_0300_),
    .B1(_0302_),
    .B2(_0308_),
    .Y(_0046_)
);

sky130_fd_sc_hd__buf_1 _1103_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[2] ),
    .X(_0309_)
);

sky130_fd_sc_hd__or2_4 _1104_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0309_),
    .B(_0302_),
    .X(_0310_)
);

sky130_fd_sc_hd__inv_8 _1105_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0310_),
    .Y(_0311_)
);

sky130_fd_sc_hd__a21o_4 _1106_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0309_),
    .A2(_0302_),
    .B1(_0311_),
    .X(_0312_)
);

sky130_fd_sc_hd__buf_1 _1107_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0145_),
    .X(_0313_)
);

sky130_fd_sc_hd__buf_1 _1108_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[2] ),
    .X(_0314_)
);

sky130_fd_sc_hd__or2_4 _1109_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0314_),
    .B(_0297_),
    .X(_0315_)
);

sky130_fd_sc_hd__inv_8 _1110_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0315_),
    .Y(_0316_)
);

sky130_fd_sc_hd__a21o_4 _1111_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0314_),
    .A2(_0297_),
    .B1(_0316_),
    .X(_0317_)
);

sky130_fd_sc_hd__o22a_4 _1112_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0272_),
    .A2(_0312_),
    .B1(_0313_),
    .B2(_0317_),
    .X(_0047_)
);

sky130_fd_sc_hd__buf_1 _1113_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0307_),
    .X(_0069_)
);

sky130_fd_sc_hd__buf_1 _1114_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[3] ),
    .X(_0318_)
);

sky130_fd_sc_hd__inv_8 _1115_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0318_),
    .Y(_0319_)
);

sky130_fd_sc_hd__buf_1 _1116_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0319_),
    .X(_0320_)
);

sky130_fd_sc_hd__or2_4 _1117_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0318_),
    .B(_0310_),
    .X(_0321_)
);

sky130_fd_sc_hd__o21a_4 _1118_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0320_),
    .A2(_0311_),
    .B1(_0321_),
    .X(_0322_)
);

sky130_fd_sc_hd__buf_1 _1119_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(P_CLK),
    .X(_0323_)
);

sky130_fd_sc_hd__inv_8 _1120_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[3] ),
    .Y(_0324_)
);

sky130_fd_sc_hd__buf_1 _1121_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0324_),
    .X(_0325_)
);

sky130_fd_sc_hd__buf_1 _1122_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[3] ),
    .X(_0326_)
);

sky130_fd_sc_hd__or2_4 _1123_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0326_),
    .B(_0315_),
    .X(_0327_)
);

sky130_fd_sc_hd__o21a_4 _1124_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0325_),
    .A2(_0316_),
    .B1(_0327_),
    .X(_0328_)
);

sky130_fd_sc_hd__a22oi_4 _1125_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0069_),
    .A2(_0322_),
    .B1(_0323_),
    .B2(_0328_),
    .Y(_0048_)
);

sky130_fd_sc_hd__buf_1 _1126_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(P_CLK),
    .X(_0329_)
);

sky130_fd_sc_hd__buf_1 _1127_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[4] ),
    .X(_0330_)
);

sky130_fd_sc_hd__or2_4 _1128_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0330_),
    .B(_0321_),
    .X(_0331_)
);

sky130_fd_sc_hd__inv_8 _1129_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0331_),
    .Y(_0332_)
);

sky130_fd_sc_hd__a21o_4 _1130_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0330_),
    .A2(_0321_),
    .B1(_0332_),
    .X(_0333_)
);

sky130_fd_sc_hd__buf_1 _1131_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[4] ),
    .X(_0334_)
);

sky130_fd_sc_hd__or2_4 _1132_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0334_),
    .B(_0327_),
    .X(_0335_)
);

sky130_fd_sc_hd__inv_8 _1133_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0335_),
    .Y(_0336_)
);

sky130_fd_sc_hd__a21o_4 _1134_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0334_),
    .A2(_0327_),
    .B1(_0336_),
    .X(_0337_)
);

sky130_fd_sc_hd__o22a_4 _1135_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0329_),
    .A2(_0333_),
    .B1(_0313_),
    .B2(_0337_),
    .X(_0049_)
);

sky130_fd_sc_hd__buf_1 _1136_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0307_),
    .X(_0338_)
);

sky130_fd_sc_hd__inv_8 _1137_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[5] ),
    .Y(_0339_)
);

sky130_fd_sc_hd__buf_1 _1138_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[5] ),
    .X(_0340_)
);

sky130_fd_sc_hd__or2_4 _1139_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0340_),
    .B(_0331_),
    .X(_0341_)
);

sky130_fd_sc_hd__o21a_4 _1140_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0339_),
    .A2(_0332_),
    .B1(_0341_),
    .X(_0342_)
);

sky130_fd_sc_hd__inv_8 _1141_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[5] ),
    .Y(_0343_)
);

sky130_fd_sc_hd__buf_1 _1142_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[5] ),
    .X(_0344_)
);

sky130_fd_sc_hd__or2_4 _1143_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0344_),
    .B(_0335_),
    .X(_0345_)
);

sky130_fd_sc_hd__o21a_4 _1144_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0343_),
    .A2(_0336_),
    .B1(_0345_),
    .X(_0346_)
);

sky130_fd_sc_hd__a22oi_4 _1145_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0338_),
    .A2(_0342_),
    .B1(_0323_),
    .B2(_0346_),
    .Y(_0050_)
);

sky130_fd_sc_hd__buf_1 _1146_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[6] ),
    .X(_0347_)
);

sky130_fd_sc_hd__or2_4 _1147_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0347_),
    .B(_0341_),
    .X(_0348_)
);

sky130_fd_sc_hd__inv_8 _1148_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0348_),
    .Y(_0349_)
);

sky130_fd_sc_hd__a21o_4 _1149_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0347_),
    .A2(_0341_),
    .B1(_0349_),
    .X(_0350_)
);

sky130_fd_sc_hd__or2_4 _1150_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[6] ),
    .B(_0345_),
    .X(_0351_)
);

sky130_fd_sc_hd__inv_8 _1151_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0351_),
    .Y(_0352_)
);

sky130_fd_sc_hd__a21o_4 _1152_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[6] ),
    .A2(_0345_),
    .B1(_0352_),
    .X(_0353_)
);

sky130_fd_sc_hd__o22a_4 _1153_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0329_),
    .A2(_0350_),
    .B1(_0313_),
    .B2(_0353_),
    .X(_0051_)
);

sky130_fd_sc_hd__inv_8 _1154_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[7] ),
    .Y(_0354_)
);

sky130_fd_sc_hd__buf_1 _1155_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0354_),
    .X(_0355_)
);

sky130_fd_sc_hd__buf_1 _1156_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0355_),
    .X(_0356_)
);

sky130_fd_sc_hd__or2_4 _1157_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[7] ),
    .B(_0348_),
    .X(_0357_)
);

sky130_fd_sc_hd__o21a_4 _1158_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0356_),
    .A2(_0349_),
    .B1(_0357_),
    .X(_0358_)
);

sky130_fd_sc_hd__inv_8 _1159_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[7] ),
    .Y(_0359_)
);

sky130_fd_sc_hd__buf_1 _1160_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0359_),
    .X(_0360_)
);

sky130_fd_sc_hd__buf_1 _1161_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0360_),
    .X(_0361_)
);

sky130_fd_sc_hd__or2_4 _1162_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[7] ),
    .B(_0351_),
    .X(_0362_)
);

sky130_fd_sc_hd__o21a_4 _1163_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0361_),
    .A2(_0352_),
    .B1(_0362_),
    .X(_0363_)
);

sky130_fd_sc_hd__a22oi_4 _1164_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0338_),
    .A2(_0358_),
    .B1(_0323_),
    .B2(_0363_),
    .Y(_0052_)
);

sky130_fd_sc_hd__buf_1 _1165_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[8] ),
    .X(_0364_)
);

sky130_fd_sc_hd__or2_4 _1166_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0364_),
    .B(_0357_),
    .X(_0365_)
);

sky130_fd_sc_hd__inv_8 _1167_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0365_),
    .Y(_0366_)
);

sky130_fd_sc_hd__a21o_4 _1168_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0364_),
    .A2(_0357_),
    .B1(_0366_),
    .X(_0367_)
);

sky130_fd_sc_hd__buf_1 _1169_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[8] ),
    .X(_0368_)
);

sky130_fd_sc_hd__or2_4 _1170_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0368_),
    .B(_0362_),
    .X(_0369_)
);

sky130_fd_sc_hd__inv_8 _1171_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0369_),
    .Y(_0370_)
);

sky130_fd_sc_hd__a21o_4 _1172_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0368_),
    .A2(_0362_),
    .B1(_0370_),
    .X(_0371_)
);

sky130_fd_sc_hd__o22a_4 _1173_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0329_),
    .A2(_0367_),
    .B1(_0313_),
    .B2(_0371_),
    .X(_0053_)
);

sky130_fd_sc_hd__inv_8 _1174_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[9] ),
    .Y(_0372_)
);

sky130_fd_sc_hd__buf_1 _1175_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0372_),
    .X(_0373_)
);

sky130_fd_sc_hd__buf_1 _1176_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0373_),
    .X(_0374_)
);

sky130_fd_sc_hd__or2_4 _1177_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[9] ),
    .B(_0365_),
    .X(_0375_)
);

sky130_fd_sc_hd__o21a_4 _1178_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0374_),
    .A2(_0366_),
    .B1(_0375_),
    .X(_0376_)
);

sky130_fd_sc_hd__inv_8 _1179_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[9] ),
    .Y(_0377_)
);

sky130_fd_sc_hd__buf_1 _1180_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0377_),
    .X(_0378_)
);

sky130_fd_sc_hd__buf_1 _1181_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0378_),
    .X(_0379_)
);

sky130_fd_sc_hd__or2_4 _1182_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[9] ),
    .B(_0369_),
    .X(_0380_)
);

sky130_fd_sc_hd__o21a_4 _1183_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0379_),
    .A2(_0370_),
    .B1(_0380_),
    .X(_0381_)
);

sky130_fd_sc_hd__a22oi_4 _1184_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0338_),
    .A2(_0376_),
    .B1(_0323_),
    .B2(_0381_),
    .Y(_0054_)
);

sky130_fd_sc_hd__inv_8 _1185_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[10] ),
    .Y(_0382_)
);

sky130_fd_sc_hd__buf_1 _1186_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0382_),
    .X(_0383_)
);

sky130_fd_sc_hd__buf_1 _1187_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0383_),
    .X(_0384_)
);

sky130_fd_sc_hd__a32o_4 _1188_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0379_),
    .A2(_0370_),
    .A3(\COUNT_BB_ONE_MIN[10] ),
    .B1(_0384_),
    .B2(_0380_),
    .X(_0385_)
);

sky130_fd_sc_hd__inv_8 _1189_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[10] ),
    .Y(_0386_)
);

sky130_fd_sc_hd__buf_1 _1190_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0386_),
    .X(_0387_)
);

sky130_fd_sc_hd__buf_1 _1191_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0387_),
    .X(_0388_)
);

sky130_fd_sc_hd__a32o_4 _1192_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0374_),
    .A2(_0366_),
    .A3(\COUNT_BB_ZERO_MIN[10] ),
    .B1(_0388_),
    .B2(_0375_),
    .X(_0389_)
);

sky130_fd_sc_hd__or2_4 _1193_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0294_),
    .B(_0389_),
    .X(_0390_)
);

sky130_fd_sc_hd__o21ai_4 _1194_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0069_),
    .A2(_0385_),
    .B1(_0390_),
    .Y(_0045_)
);

sky130_fd_sc_hd__inv_8 _1195_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ZERO),
    .Y(_0391_)
);

sky130_fd_sc_hd__buf_1 _1196_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0391_),
    .X(_0392_)
);

sky130_fd_sc_hd__buf_1 _1197_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[9] ),
    .X(_0393_)
);

sky130_fd_sc_hd__buf_1 _1198_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[6] ),
    .X(_0394_)
);

sky130_fd_sc_hd__and2_4 _1199_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0355_),
    .B(_0394_),
    .X(_0395_)
);

sky130_fd_sc_hd__inv_8 _1200_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[8] ),
    .Y(_0396_)
);

sky130_fd_sc_hd__buf_1 _1201_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[7] ),
    .X(_0397_)
);

sky130_fd_sc_hd__inv_8 _1202_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[6] ),
    .Y(_0398_)
);

sky130_fd_sc_hd__buf_1 _1203_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0398_),
    .X(_0399_)
);

sky130_fd_sc_hd__buf_1 _1204_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[5] ),
    .X(_0400_)
);

sky130_fd_sc_hd__a2bb2o_4 _1205_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0396_),
    .A2_N(_0397_),
    .B1(_0399_),
    .B2(_0400_),
    .X(_0401_)
);

sky130_fd_sc_hd__inv_8 _1206_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[7] ),
    .Y(_0402_)
);

sky130_fd_sc_hd__buf_1 _1207_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0402_),
    .X(_0403_)
);

sky130_fd_sc_hd__or2_4 _1208_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0364_),
    .B(_0403_),
    .X(_0404_)
);

sky130_fd_sc_hd__o21ai_4 _1209_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0355_),
    .A2(_0394_),
    .B1(_0404_),
    .Y(_0405_)
);

sky130_fd_sc_hd__inv_8 _1210_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0400_),
    .Y(_0406_)
);

sky130_fd_sc_hd__inv_8 _1211_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[4] ),
    .Y(_0407_)
);

sky130_fd_sc_hd__buf_1 _1212_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0407_),
    .X(_0408_)
);

sky130_fd_sc_hd__or2_4 _1213_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0340_),
    .B(_0408_),
    .X(_0409_)
);

sky130_fd_sc_hd__inv_8 _1214_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[3] ),
    .Y(_0410_)
);

sky130_fd_sc_hd__buf_1 _1215_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0410_),
    .X(_0411_)
);

sky130_fd_sc_hd__inv_8 _1216_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[2] ),
    .Y(_0412_)
);

sky130_fd_sc_hd__inv_8 _1217_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[1] ),
    .Y(_0413_)
);

sky130_fd_sc_hd__inv_8 _1218_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[0] ),
    .Y(_0414_)
);

sky130_fd_sc_hd__buf_1 _1219_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0414_),
    .X(_0415_)
);

sky130_fd_sc_hd__o22a_4 _1220_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0309_),
    .A2(_0413_),
    .B1(_0301_),
    .B2(_0415_),
    .X(_0416_)
);

sky130_fd_sc_hd__and2_4 _1221_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0309_),
    .B(_0413_),
    .X(_0417_)
);

sky130_fd_sc_hd__o22a_4 _1222_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0318_),
    .A2(_0412_),
    .B1(_0416_),
    .B2(_0417_),
    .X(_0418_)
);

sky130_fd_sc_hd__buf_1 _1223_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[2] ),
    .X(_0419_)
);

sky130_fd_sc_hd__a2bb2o_4 _1224_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0319_),
    .A2_N(_0419_),
    .B1(_0330_),
    .B2(_0410_),
    .X(_0420_)
);

sky130_fd_sc_hd__o22a_4 _1225_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0330_),
    .A2(_0411_),
    .B1(_0418_),
    .B2(_0420_),
    .X(_0421_)
);

sky130_fd_sc_hd__a21o_4 _1226_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0340_),
    .A2(_0408_),
    .B1(_0421_),
    .X(_0422_)
);

sky130_fd_sc_hd__a22oi_4 _1227_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0347_),
    .A2(_0406_),
    .B1(_0409_),
    .B2(_0422_),
    .Y(_0423_)
);

sky130_fd_sc_hd__inv_8 _1228_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[6] ),
    .Y(_0424_)
);

sky130_fd_sc_hd__buf_1 _1229_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0424_),
    .X(_0425_)
);

sky130_fd_sc_hd__a32oi_4 _1230_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO_MIN[7] ),
    .A2(_0425_),
    .A3(_0404_),
    .B1(_0364_),
    .B2(_0403_),
    .Y(_0426_)
);

sky130_fd_sc_hd__o41a_4 _1231_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0395_),
    .A2(_0401_),
    .A3(_0405_),
    .A4(_0423_),
    .B1(_0426_),
    .X(_0427_)
);

sky130_fd_sc_hd__buf_1 _1232_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[8] ),
    .X(_0428_)
);

sky130_fd_sc_hd__a2bb2o_4 _1233_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0387_),
    .A2_N(_0393_),
    .B1(_0373_),
    .B2(_0428_),
    .X(_0429_)
);

sky130_fd_sc_hd__o22a_4 _1234_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0386_),
    .A2(_0393_),
    .B1(_0373_),
    .B2(_0428_),
    .X(_0430_)
);

sky130_fd_sc_hd__o21a_4 _1235_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0427_),
    .A2(_0429_),
    .B1(_0430_),
    .X(_0431_)
);

sky130_fd_sc_hd__a211o_4 _1236_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0387_),
    .A2(_0393_),
    .B1(\COUNT_BB_ZERO[10] ),
    .C1(_0431_),
    .X(_0432_)
);

sky130_fd_sc_hd__inv_8 _1237_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0432_),
    .Y(_0433_)
);

sky130_fd_sc_hd__or4_4 _1238_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[8] ),
    .B(\COUNT_BB_ZERO[7] ),
    .C(\COUNT_BB_ZERO[6] ),
    .D(\COUNT_BB_ZERO[5] ),
    .X(_0434_)
);

sky130_fd_sc_hd__or4_4 _1239_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[4] ),
    .B(\COUNT_BB_ZERO[3] ),
    .C(\COUNT_BB_ZERO[2] ),
    .D(\COUNT_BB_ZERO[1] ),
    .X(_0435_)
);

sky130_fd_sc_hd__nor4_4 _1240_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[10] ),
    .B(\COUNT_BB_ZERO[9] ),
    .C(_0434_),
    .D(_0435_),
    .Y(_0436_)
);

sky130_fd_sc_hd__and2_4 _1241_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0433_),
    .B(_0436_),
    .X(_0437_)
);

sky130_fd_sc_hd__or2_4 _1242_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0306_),
    .B(_0437_),
    .X(_0438_)
);

sky130_fd_sc_hd__buf_1 _1243_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0438_),
    .X(_0439_)
);

sky130_fd_sc_hd__inv_8 _1244_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0439_),
    .Y(_0440_)
);

sky130_fd_sc_hd__and2_4 _1245_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0306_),
    .B(_0437_),
    .X(_0441_)
);

sky130_fd_sc_hd__inv_8 _1246_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[10] ),
    .Y(_0442_)
);

sky130_fd_sc_hd__buf_1 _1247_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0442_),
    .X(_0443_)
);

sky130_fd_sc_hd__inv_8 _1248_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[9]),
    .Y(_0444_)
);

sky130_fd_sc_hd__and2_4 _1249_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0372_),
    .B(_0444_),
    .X(_0445_)
);

sky130_fd_sc_hd__buf_1 _1250_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0396_),
    .X(_0446_)
);

sky130_fd_sc_hd__inv_8 _1251_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[8]),
    .Y(_0447_)
);

sky130_fd_sc_hd__and2_4 _1252_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0396_),
    .B(_0447_),
    .X(_0448_)
);

sky130_fd_sc_hd__inv_8 _1253_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[7]),
    .Y(_0449_)
);

sky130_fd_sc_hd__and2_4 _1254_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0354_),
    .B(_0449_),
    .X(_0450_)
);

sky130_fd_sc_hd__inv_8 _1255_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[6]),
    .Y(_0451_)
);

sky130_fd_sc_hd__buf_1 _1256_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0451_),
    .X(_0452_)
);

sky130_fd_sc_hd__a2bb2o_4 _1257_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0398_),
    .A2_N(_0452_),
    .B1(_0398_),
    .B2(_0451_),
    .X(_0453_)
);

sky130_fd_sc_hd__inv_8 _1258_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[5]),
    .Y(_0454_)
);

sky130_fd_sc_hd__or2_4 _1259_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[5] ),
    .B(SCAN_IN[5]),
    .X(_0455_)
);

sky130_fd_sc_hd__o21ai_4 _1260_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0339_),
    .A2(_0454_),
    .B1(_0455_),
    .Y(_0456_)
);

sky130_fd_sc_hd__inv_8 _1261_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[4] ),
    .Y(_0457_)
);

sky130_fd_sc_hd__inv_8 _1262_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[4]),
    .Y(_0458_)
);

sky130_fd_sc_hd__buf_1 _1263_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0458_),
    .X(_0459_)
);

sky130_fd_sc_hd__a2bb2o_4 _1264_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0457_),
    .A2_N(_0459_),
    .B1(_0457_),
    .B2(_0458_),
    .X(_0460_)
);

sky130_fd_sc_hd__inv_8 _1265_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[3]),
    .Y(_0461_)
);

sky130_fd_sc_hd__or2_4 _1266_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[3] ),
    .B(SCAN_IN[3]),
    .X(_0462_)
);

sky130_fd_sc_hd__o21ai_4 _1267_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0319_),
    .A2(_0461_),
    .B1(_0462_),
    .Y(_0463_)
);

sky130_fd_sc_hd__inv_8 _1268_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[2] ),
    .Y(_0464_)
);

sky130_fd_sc_hd__inv_8 _1269_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[2]),
    .Y(_0465_)
);

sky130_fd_sc_hd__a2bb2o_4 _1270_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0464_),
    .A2_N(_0465_),
    .B1(_0464_),
    .B2(_0465_),
    .X(_0466_)
);

sky130_fd_sc_hd__and2_4 _1271_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[0] ),
    .B(SCAN_IN[0]),
    .X(_0467_)
);

sky130_fd_sc_hd__inv_8 _1272_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[1]),
    .Y(_0468_)
);

sky130_fd_sc_hd__o22a_4 _1273_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0303_),
    .A2(_0468_),
    .B1(_0301_),
    .B2(SCAN_IN[1]),
    .X(_0469_)
);

sky130_fd_sc_hd__and2_4 _1274_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0467_),
    .B(_0469_),
    .X(_0470_)
);

sky130_fd_sc_hd__a21oi_4 _1275_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0301_),
    .A2(SCAN_IN[1]),
    .B1(_0470_),
    .Y(_0471_)
);

sky130_fd_sc_hd__nor3_4 _1276_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0463_),
    .B(_0466_),
    .C(_0471_),
    .Y(_0472_)
);

sky130_fd_sc_hd__a32o_4 _1277_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO_MIN[2] ),
    .A2(SCAN_IN[2]),
    .A3(_0462_),
    .B1(_0318_),
    .B2(SCAN_IN[3]),
    .X(_0473_)
);

sky130_fd_sc_hd__nor2_4 _1278_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0472_),
    .B(_0473_),
    .Y(_0474_)
);

sky130_fd_sc_hd__nor3_4 _1279_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0456_),
    .B(_0460_),
    .C(_0474_),
    .Y(_0475_)
);

sky130_fd_sc_hd__a32o_4 _1280_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0330_),
    .A2(SCAN_IN[4]),
    .A3(_0455_),
    .B1(\COUNT_BB_ZERO_MIN[5] ),
    .B2(SCAN_IN[5]),
    .X(_0476_)
);

sky130_fd_sc_hd__nor2_4 _1281_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0475_),
    .B(_0476_),
    .Y(_0477_)
);

sky130_fd_sc_hd__o22a_4 _1282_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0398_),
    .A2(_0452_),
    .B1(_0453_),
    .B2(_0477_),
    .X(_0478_)
);

sky130_fd_sc_hd__o22a_4 _1283_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0355_),
    .A2(_0449_),
    .B1(_0450_),
    .B2(_0478_),
    .X(_0479_)
);

sky130_fd_sc_hd__o22a_4 _1284_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0446_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0479_),
    .X(_0480_)
);

sky130_fd_sc_hd__o22a_4 _1285_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0373_),
    .A2(_0444_),
    .B1(_0445_),
    .B2(_0480_),
    .X(_0481_)
);

sky130_fd_sc_hd__inv_8 _1286_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[10]),
    .Y(_0482_)
);

sky130_fd_sc_hd__o22a_4 _1287_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0387_),
    .A2(SCAN_IN[10]),
    .B1(\COUNT_BB_ZERO_MIN[10] ),
    .B2(_0482_),
    .X(_0483_)
);

sky130_fd_sc_hd__xor2_4 _1288_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0481_),
    .B(_0483_),
    .X(_0484_)
);

sky130_fd_sc_hd__buf_1 _1289_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0393_),
    .X(_0485_)
);

sky130_fd_sc_hd__a21oi_4 _1290_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO_MIN[8] ),
    .A2(SCAN_IN[8]),
    .B1(_0448_),
    .Y(_0486_)
);

sky130_fd_sc_hd__xor2_4 _1291_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0479_),
    .B(_0486_),
    .X(_0487_)
);

sky130_fd_sc_hd__a21o_4 _1292_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO_MIN[7] ),
    .A2(SCAN_IN[7]),
    .B1(_0450_),
    .X(_0488_)
);

sky130_fd_sc_hd__a2bb2o_4 _1293_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0478_),
    .A2_N(_0488_),
    .B1(_0478_),
    .B2(_0488_),
    .X(_0489_)
);

sky130_fd_sc_hd__and2_4 _1294_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[7] ),
    .B(_0489_),
    .X(_0490_)
);

sky130_fd_sc_hd__a2bb2oi_4 _1295_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0453_),
    .A2_N(_0477_),
    .B1(_0453_),
    .B2(_0477_),
    .Y(_0491_)
);

sky130_fd_sc_hd__nor2_4 _1296_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0424_),
    .B(_0491_),
    .Y(_0492_)
);

sky130_fd_sc_hd__and2_4 _1297_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0424_),
    .B(_0491_),
    .X(_0493_)
);

sky130_fd_sc_hd__o22a_4 _1298_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0457_),
    .A2(_0459_),
    .B1(_0474_),
    .B2(_0460_),
    .X(_0494_)
);

sky130_fd_sc_hd__a2bb2o_4 _1299_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0456_),
    .A2_N(_0494_),
    .B1(_0456_),
    .B2(_0494_),
    .X(_0495_)
);

sky130_fd_sc_hd__nor2_4 _1300_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[5] ),
    .B(_0495_),
    .Y(_0496_)
);

sky130_fd_sc_hd__and2_4 _1301_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[5] ),
    .B(_0495_),
    .X(_0497_)
);

sky130_fd_sc_hd__a2bb2oi_4 _1302_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0474_),
    .A2_N(_0460_),
    .B1(_0474_),
    .B2(_0460_),
    .Y(_0498_)
);

sky130_fd_sc_hd__nor2_4 _1303_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0408_),
    .B(_0498_),
    .Y(_0499_)
);

sky130_fd_sc_hd__buf_1 _1304_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0464_),
    .X(_0500_)
);

sky130_fd_sc_hd__o22a_4 _1305_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0500_),
    .A2(_0465_),
    .B1(_0471_),
    .B2(_0466_),
    .X(_0501_)
);

sky130_fd_sc_hd__a2bb2oi_4 _1306_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0463_),
    .A2_N(_0501_),
    .B1(_0463_),
    .B2(_0501_),
    .Y(_0502_)
);

sky130_fd_sc_hd__and2_4 _1307_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0411_),
    .B(_0502_),
    .X(_0503_)
);

sky130_fd_sc_hd__and2_4 _1308_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0407_),
    .B(_0498_),
    .X(_0504_)
);

sky130_fd_sc_hd__a2bb2o_4 _1309_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0471_),
    .A2_N(_0466_),
    .B1(_0471_),
    .B2(_0466_),
    .X(_0505_)
);

sky130_fd_sc_hd__inv_8 _1310_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0469_),
    .Y(_0506_)
);

sky130_fd_sc_hd__or2_4 _1311_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[0] ),
    .B(SCAN_IN[0]),
    .X(_0507_)
);

sky130_fd_sc_hd__a21o_4 _1312_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0414_),
    .A2(_0507_),
    .B1(_0467_),
    .X(_0508_)
);

sky130_fd_sc_hd__a21oi_4 _1313_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0413_),
    .A2(_0469_),
    .B1(_0508_),
    .Y(_0509_)
);

sky130_fd_sc_hd__a211o_4 _1314_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO[1] ),
    .A2(_0506_),
    .B1(_0470_),
    .C1(_0509_),
    .X(_0510_)
);

sky130_fd_sc_hd__a21oi_4 _1315_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0505_),
    .A2(_0510_),
    .B1(\COUNT_BB_ZERO[2] ),
    .Y(_0511_)
);

sky130_fd_sc_hd__nor2_4 _1316_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0505_),
    .B(_0510_),
    .Y(_0512_)
);

sky130_fd_sc_hd__o22a_4 _1317_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0411_),
    .A2(_0502_),
    .B1(_0511_),
    .B2(_0512_),
    .X(_0513_)
);

sky130_fd_sc_hd__nor3_4 _1318_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0503_),
    .B(_0504_),
    .C(_0513_),
    .Y(_0514_)
);

sky130_fd_sc_hd__nor3_4 _1319_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0497_),
    .B(_0499_),
    .C(_0514_),
    .Y(_0515_)
);

sky130_fd_sc_hd__nor3_4 _1320_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0493_),
    .B(_0496_),
    .C(_0515_),
    .Y(_0516_)
);

sky130_fd_sc_hd__nor3_4 _1321_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0490_),
    .B(_0492_),
    .C(_0516_),
    .Y(_0517_)
);

sky130_fd_sc_hd__or2_4 _1322_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0397_),
    .B(_0489_),
    .X(_0518_)
);

sky130_fd_sc_hd__o21ai_4 _1323_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO[8] ),
    .A2(_0487_),
    .B1(_0518_),
    .Y(_0519_)
);

sky130_fd_sc_hd__or2_4 _1324_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0517_),
    .B(_0519_),
    .X(_0520_)
);

sky130_fd_sc_hd__a21bo_4 _1325_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0428_),
    .A2(_0487_),
    .B1_N(_0520_),
    .X(_0521_)
);

sky130_fd_sc_hd__nor2_4 _1326_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0485_),
    .B(_0521_),
    .Y(_0522_)
);

sky130_fd_sc_hd__a21o_4 _1327_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO_MIN[9] ),
    .A2(SCAN_IN[9]),
    .B1(_0445_),
    .X(_0523_)
);

sky130_fd_sc_hd__a2bb2oi_4 _1328_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0480_),
    .A2_N(_0523_),
    .B1(_0480_),
    .B2(_0523_),
    .Y(_0524_)
);

sky130_fd_sc_hd__a21boi_4 _1329_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0485_),
    .A2(_0521_),
    .B1_N(_0524_),
    .Y(_0525_)
);

sky130_fd_sc_hd__a211o_4 _1330_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0442_),
    .A2(_0484_),
    .B1(_0522_),
    .C1(_0525_),
    .X(_0526_)
);

sky130_fd_sc_hd__o21ai_4 _1331_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0443_),
    .A2(_0484_),
    .B1(_0526_),
    .Y(_0527_)
);

sky130_fd_sc_hd__inv_8 _1332_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0393_),
    .Y(_0528_)
);

sky130_fd_sc_hd__or2_4 _1333_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0528_),
    .B(SCAN_IN[20]),
    .X(_0529_)
);

sky130_fd_sc_hd__buf_1 _1334_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[1] ),
    .X(_0530_)
);

sky130_fd_sc_hd__inv_8 _1335_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[12]),
    .Y(_0531_)
);

sky130_fd_sc_hd__and2_4 _1336_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0413_),
    .B(SCAN_IN[12]),
    .X(_0532_)
);

sky130_fd_sc_hd__nor2_4 _1337_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[11]),
    .B(_0415_),
    .Y(_0533_)
);

sky130_fd_sc_hd__a211o_4 _1338_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0530_),
    .A2(_0531_),
    .B1(_0532_),
    .C1(_0533_),
    .X(_0534_)
);

sky130_fd_sc_hd__inv_8 _1339_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[13]),
    .Y(_0535_)
);

sky130_fd_sc_hd__buf_1 _1340_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[3] ),
    .X(_0536_)
);

sky130_fd_sc_hd__inv_8 _1341_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[14]),
    .Y(_0537_)
);

sky130_fd_sc_hd__and2_4 _1342_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0536_),
    .B(_0537_),
    .X(_0538_)
);

sky130_fd_sc_hd__o22a_4 _1343_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0536_),
    .A2(_0537_),
    .B1(_0419_),
    .B2(_0535_),
    .X(_0539_)
);

sky130_fd_sc_hd__inv_8 _1344_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0539_),
    .Y(_0540_)
);

sky130_fd_sc_hd__a211o_4 _1345_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0419_),
    .A2(_0535_),
    .B1(_0538_),
    .C1(_0540_),
    .X(_0541_)
);

sky130_fd_sc_hd__inv_8 _1346_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[20]),
    .Y(_0542_)
);

sky130_fd_sc_hd__inv_8 _1347_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[15]),
    .Y(_0543_)
);

sky130_fd_sc_hd__buf_1 _1348_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[4] ),
    .X(_0544_)
);

sky130_fd_sc_hd__and2_4 _1349_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0543_),
    .B(_0544_),
    .X(_0545_)
);

sky130_fd_sc_hd__and2_4 _1350_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[11]),
    .B(_0415_),
    .X(_0546_)
);

sky130_fd_sc_hd__inv_8 _1351_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[17]),
    .Y(_0547_)
);

sky130_fd_sc_hd__or2_4 _1352_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0402_),
    .B(SCAN_IN[18]),
    .X(_0548_)
);

sky130_fd_sc_hd__buf_1 _1353_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0548_),
    .X(_0549_)
);

sky130_fd_sc_hd__inv_8 _1354_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0549_),
    .Y(_0550_)
);

sky130_fd_sc_hd__a2bb2o_4 _1355_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(\COUNT_BB_ZERO[6] ),
    .A2_N(_0547_),
    .B1(_0402_),
    .B2(SCAN_IN[18]),
    .X(_0551_)
);

sky130_fd_sc_hd__a211o_4 _1356_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0394_),
    .A2(_0547_),
    .B1(_0550_),
    .C1(_0551_),
    .X(_0552_)
);

sky130_fd_sc_hd__a2111o_4 _1357_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO[9] ),
    .A2(_0542_),
    .B1(_0545_),
    .C1(_0546_),
    .D1(_0552_),
    .X(_0553_)
);

sky130_fd_sc_hd__inv_8 _1358_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[8] ),
    .Y(_0554_)
);

sky130_fd_sc_hd__or2_4 _1359_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0554_),
    .B(SCAN_IN[19]),
    .X(_0555_)
);

sky130_fd_sc_hd__buf_1 _1360_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0555_),
    .X(_0556_)
);

sky130_fd_sc_hd__or2_4 _1361_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0406_),
    .B(SCAN_IN[16]),
    .X(_0557_)
);

sky130_fd_sc_hd__inv_8 _1362_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[19]),
    .Y(_0558_)
);

sky130_fd_sc_hd__o22a_4 _1363_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ZERO[8] ),
    .A2(_0558_),
    .B1(\COUNT_BB_ZERO[9] ),
    .B2(_0542_),
    .X(_0559_)
);

sky130_fd_sc_hd__inv_8 _1364_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[16]),
    .Y(_0560_)
);

sky130_fd_sc_hd__o22a_4 _1365_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0400_),
    .A2(_0560_),
    .B1(_0543_),
    .B2(_0544_),
    .X(_0561_)
);

sky130_fd_sc_hd__nand4_4 _1366_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0556_),
    .B(_0557_),
    .C(_0559_),
    .D(_0561_),
    .Y(_0562_)
);

sky130_fd_sc_hd__or4_4 _1367_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0534_),
    .B(_0541_),
    .C(_0553_),
    .D(_0562_),
    .X(_0563_)
);

sky130_fd_sc_hd__inv_8 _1368_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0556_),
    .Y(_0564_)
);

sky130_fd_sc_hd__inv_8 _1369_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0552_),
    .Y(_0565_)
);

sky130_fd_sc_hd__o21a_4 _1370_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0530_),
    .A2(_0531_),
    .B1(_0534_),
    .X(_0566_)
);

sky130_fd_sc_hd__o22a_4 _1371_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0566_),
    .A2(_0541_),
    .B1(_0539_),
    .B2(_0538_),
    .X(_0567_)
);

sky130_fd_sc_hd__o21ai_4 _1372_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0545_),
    .A2(_0567_),
    .B1(_0561_),
    .Y(_0568_)
);

sky130_fd_sc_hd__a32oi_4 _1373_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0565_),
    .A2(_0557_),
    .A3(_0568_),
    .B1(_0551_),
    .B2(_0549_),
    .Y(_0569_)
);

sky130_fd_sc_hd__o21ai_4 _1374_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0564_),
    .A2(_0569_),
    .B1(_0559_),
    .Y(_0570_)
);

sky130_fd_sc_hd__a32o_4 _1375_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0529_),
    .A2(_0563_),
    .A3(_0570_),
    .B1(SCAN_IN[21]),
    .B2(_0442_),
    .X(_0571_)
);

sky130_fd_sc_hd__o21a_4 _1376_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[21]),
    .A2(_0443_),
    .B1(_0571_),
    .X(_0572_)
);

sky130_fd_sc_hd__or2_4 _1377_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0527_),
    .B(_0572_),
    .X(_0573_)
);

sky130_fd_sc_hd__buf_1 _1378_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0573_),
    .X(_0574_)
);

sky130_fd_sc_hd__and2_4 _1379_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0306_),
    .B(_0574_),
    .X(_0575_)
);

sky130_fd_sc_hd__buf_1 _1380_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ZERO),
    .X(_0576_)
);

sky130_fd_sc_hd__buf_1 _1381_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0572_),
    .X(_0577_)
);

sky130_fd_sc_hd__buf_1 _1382_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0527_),
    .X(_0578_)
);

sky130_fd_sc_hd__nor3_4 _1383_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO[0] ),
    .B(_0577_),
    .C(_0578_),
    .Y(_0579_)
);

sky130_fd_sc_hd__or2_4 _1384_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0576_),
    .B(_0579_),
    .X(_0580_)
);

sky130_fd_sc_hd__o32ai_4 _1385_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0392_),
    .A2(_0440_),
    .A3(_0441_),
    .B1(_0575_),
    .B2(_0580_),
    .Y(_0034_)
);

sky130_fd_sc_hd__or3_4 _1386_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0530_),
    .B(_0577_),
    .C(_0578_),
    .X(_0581_)
);

sky130_fd_sc_hd__nand2_4 _1387_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0304_),
    .B(_0574_),
    .Y(_0582_)
);

sky130_fd_sc_hd__buf_1 _1388_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0433_),
    .X(_0583_)
);

sky130_fd_sc_hd__o22a_4 _1389_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0301_),
    .A2(_0583_),
    .B1(_0304_),
    .B2(_0432_),
    .X(_0584_)
);

sky130_fd_sc_hd__nand2_4 _1390_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0439_),
    .B(_0584_),
    .Y(_0585_)
);

sky130_fd_sc_hd__o21a_4 _1391_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0439_),
    .A2(_0584_),
    .B1(_0576_),
    .X(_0586_)
);

sky130_fd_sc_hd__a32o_4 _1392_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0392_),
    .A2(_0581_),
    .A3(_0582_),
    .B1(_0585_),
    .B2(_0586_),
    .X(_0036_)
);

sky130_fd_sc_hd__and2_4 _1393_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0500_),
    .B(_0574_),
    .X(_0587_)
);

sky130_fd_sc_hd__nor3_4 _1394_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0419_),
    .B(_0577_),
    .C(_0578_),
    .Y(_0588_)
);

sky130_fd_sc_hd__or2_4 _1395_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0576_),
    .B(_0588_),
    .X(_0589_)
);

sky130_fd_sc_hd__buf_1 _1396_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0432_),
    .X(_0590_)
);

sky130_fd_sc_hd__or3_4 _1397_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0303_),
    .B(_0305_),
    .C(_0436_),
    .X(_0591_)
);

sky130_fd_sc_hd__or2_4 _1398_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0500_),
    .B(_0591_),
    .X(_0592_)
);

sky130_fd_sc_hd__inv_8 _1399_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0592_),
    .Y(_0593_)
);

sky130_fd_sc_hd__a21oi_4 _1400_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0500_),
    .A2(_0591_),
    .B1(_0593_),
    .Y(_0594_)
);

sky130_fd_sc_hd__or2_4 _1401_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0590_),
    .B(_0594_),
    .X(_0595_)
);

sky130_fd_sc_hd__buf_1 _1402_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ZERO),
    .X(_0596_)
);

sky130_fd_sc_hd__o21a_4 _1403_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0312_),
    .A2(_0583_),
    .B1(_0596_),
    .X(_0597_)
);

sky130_fd_sc_hd__a2bb2o_4 _1404_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0587_),
    .A2_N(_0589_),
    .B1(_0595_),
    .B2(_0597_),
    .X(_0037_)
);

sky130_fd_sc_hd__buf_1 _1405_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0576_),
    .X(_0598_)
);

sky130_fd_sc_hd__buf_1 _1406_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0572_),
    .X(_0599_)
);

sky130_fd_sc_hd__buf_1 _1407_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0527_),
    .X(_0600_)
);

sky130_fd_sc_hd__nor3_4 _1408_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0536_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0601_)
);

sky130_fd_sc_hd__and2_4 _1409_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0320_),
    .B(_0574_),
    .X(_0602_)
);

sky130_fd_sc_hd__or2_4 _1410_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0318_),
    .B(_0593_),
    .X(_0603_)
);

sky130_fd_sc_hd__or2_4 _1411_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0320_),
    .B(_0592_),
    .X(_0604_)
);

sky130_fd_sc_hd__buf_1 _1412_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0432_),
    .X(_0605_)
);

sky130_fd_sc_hd__a21oi_4 _1413_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0603_),
    .A2(_0604_),
    .B1(_0605_),
    .Y(_0606_)
);

sky130_fd_sc_hd__a21o_4 _1414_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0322_),
    .A2(_0605_),
    .B1(_0392_),
    .X(_0607_)
);

sky130_fd_sc_hd__o32ai_4 _1415_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0598_),
    .A2(_0601_),
    .A3(_0602_),
    .B1(_0606_),
    .B2(_0607_),
    .Y(_0038_)
);

sky130_fd_sc_hd__nor3_4 _1416_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0544_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0608_)
);

sky130_fd_sc_hd__buf_1 _1417_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0457_),
    .X(_0609_)
);

sky130_fd_sc_hd__buf_1 _1418_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0573_),
    .X(_0610_)
);

sky130_fd_sc_hd__and2_4 _1419_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0609_),
    .B(_0610_),
    .X(_0611_)
);

sky130_fd_sc_hd__buf_1 _1420_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0583_),
    .X(_0612_)
);

sky130_fd_sc_hd__nor2_4 _1421_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0333_),
    .B(_0612_),
    .Y(_0613_)
);

sky130_fd_sc_hd__or2_4 _1422_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0609_),
    .B(_0604_),
    .X(_0614_)
);

sky130_fd_sc_hd__inv_8 _1423_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0614_),
    .Y(_0615_)
);

sky130_fd_sc_hd__a21o_4 _1424_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0609_),
    .A2(_0604_),
    .B1(_0615_),
    .X(_0616_)
);

sky130_fd_sc_hd__a21o_4 _1425_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0612_),
    .A2(_0616_),
    .B1(_0392_),
    .X(_0617_)
);

sky130_fd_sc_hd__o32ai_4 _1426_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0598_),
    .A2(_0608_),
    .A3(_0611_),
    .B1(_0613_),
    .B2(_0617_),
    .Y(_0039_)
);

sky130_fd_sc_hd__nor3_4 _1427_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0400_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0618_)
);

sky130_fd_sc_hd__and2_4 _1428_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0339_),
    .B(_0610_),
    .X(_0619_)
);

sky130_fd_sc_hd__or2_4 _1429_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0340_),
    .B(_0615_),
    .X(_0620_)
);

sky130_fd_sc_hd__or2_4 _1430_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0339_),
    .B(_0614_),
    .X(_0621_)
);

sky130_fd_sc_hd__a21oi_4 _1431_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0620_),
    .A2(_0621_),
    .B1(_0605_),
    .Y(_0622_)
);

sky130_fd_sc_hd__a21o_4 _1432_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0342_),
    .A2(_0605_),
    .B1(_0392_),
    .X(_0623_)
);

sky130_fd_sc_hd__o32ai_4 _1433_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0598_),
    .A2(_0618_),
    .A3(_0619_),
    .B1(_0622_),
    .B2(_0623_),
    .Y(_0040_)
);

sky130_fd_sc_hd__and2_4 _1434_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0399_),
    .B(_0574_),
    .X(_0624_)
);

sky130_fd_sc_hd__nor3_4 _1435_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0394_),
    .B(_0577_),
    .C(_0578_),
    .Y(_0625_)
);

sky130_fd_sc_hd__or2_4 _1436_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0576_),
    .B(_0625_),
    .X(_0626_)
);

sky130_fd_sc_hd__or2_4 _1437_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0399_),
    .B(_0621_),
    .X(_0627_)
);

sky130_fd_sc_hd__a21boi_4 _1438_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0399_),
    .A2(_0621_),
    .B1_N(_0627_),
    .Y(_0628_)
);

sky130_fd_sc_hd__or2_4 _1439_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0590_),
    .B(_0628_),
    .X(_0629_)
);

sky130_fd_sc_hd__o21a_4 _1440_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0350_),
    .A2(_0583_),
    .B1(_0596_),
    .X(_0630_)
);

sky130_fd_sc_hd__a2bb2o_4 _1441_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0624_),
    .A2_N(_0626_),
    .B1(_0629_),
    .B2(_0630_),
    .X(_0041_)
);

sky130_fd_sc_hd__nor3_4 _1442_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0397_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0631_)
);

sky130_fd_sc_hd__and2_4 _1443_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0356_),
    .B(_0610_),
    .X(_0632_)
);

sky130_fd_sc_hd__and2_4 _1444_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0356_),
    .B(_0627_),
    .X(_0633_)
);

sky130_fd_sc_hd__or2_4 _1445_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0356_),
    .B(_0627_),
    .X(_0634_)
);

sky130_fd_sc_hd__buf_1 _1446_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0634_),
    .X(_0635_)
);

sky130_fd_sc_hd__inv_8 _1447_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0635_),
    .Y(_0636_)
);

sky130_fd_sc_hd__o21a_4 _1448_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0633_),
    .A2(_0636_),
    .B1(_0612_),
    .X(_0637_)
);

sky130_fd_sc_hd__a21o_4 _1449_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0358_),
    .A2(_0590_),
    .B1(_0391_),
    .X(_0638_)
);

sky130_fd_sc_hd__o32ai_4 _1450_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0598_),
    .A2(_0631_),
    .A3(_0632_),
    .B1(_0637_),
    .B2(_0638_),
    .Y(_0042_)
);

sky130_fd_sc_hd__nor3_4 _1451_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0428_),
    .B(_0577_),
    .C(_0578_),
    .Y(_0639_)
);

sky130_fd_sc_hd__and2_4 _1452_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0446_),
    .B(_0573_),
    .X(_0640_)
);

sky130_fd_sc_hd__nor3_4 _1453_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0596_),
    .B(_0639_),
    .C(_0640_),
    .Y(_0641_)
);

sky130_fd_sc_hd__or2_4 _1454_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0446_),
    .B(_0635_),
    .X(_0642_)
);

sky130_fd_sc_hd__inv_8 _1455_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0642_),
    .Y(_0643_)
);

sky130_fd_sc_hd__a21o_4 _1456_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0446_),
    .A2(_0635_),
    .B1(_0643_),
    .X(_0644_)
);

sky130_fd_sc_hd__o21a_4 _1457_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0367_),
    .A2(_0583_),
    .B1(MULTIBIT_ZERO),
    .X(_0645_)
);

sky130_fd_sc_hd__a21boi_4 _1458_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0612_),
    .A2(_0644_),
    .B1_N(_0645_),
    .Y(_0646_)
);

sky130_fd_sc_hd__or2_4 _1459_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0641_),
    .B(_0646_),
    .X(_0043_)
);

sky130_fd_sc_hd__nor3_4 _1460_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0485_),
    .B(_0599_),
    .C(_0600_),
    .Y(_0647_)
);

sky130_fd_sc_hd__and2_4 _1461_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0374_),
    .B(_0610_),
    .X(_0648_)
);

sky130_fd_sc_hd__and2_4 _1462_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0374_),
    .B(_0642_),
    .X(_0649_)
);

sky130_fd_sc_hd__and2_4 _1463_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ZERO_MIN[9] ),
    .B(_0643_),
    .X(_0650_)
);

sky130_fd_sc_hd__o21a_4 _1464_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0649_),
    .A2(_0650_),
    .B1(_0612_),
    .X(_0651_)
);

sky130_fd_sc_hd__a21o_4 _1465_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0376_),
    .A2(_0590_),
    .B1(_0391_),
    .X(_0652_)
);

sky130_fd_sc_hd__o32ai_4 _1466_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0596_),
    .A2(_0647_),
    .A3(_0648_),
    .B1(_0651_),
    .B2(_0652_),
    .Y(_0044_)
);

sky130_fd_sc_hd__inv_8 _1467_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0571_),
    .Y(_0653_)
);

sky130_fd_sc_hd__and3_4 _1468_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0443_),
    .B(_0653_),
    .C(_0526_),
    .X(_0654_)
);

sky130_fd_sc_hd__and2_4 _1469_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0388_),
    .B(_0610_),
    .X(_0655_)
);

sky130_fd_sc_hd__and2_4 _1470_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0388_),
    .B(_0650_),
    .X(_0656_)
);

sky130_fd_sc_hd__nor2_4 _1471_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0388_),
    .B(_0650_),
    .Y(_0657_)
);

sky130_fd_sc_hd__nor3_4 _1472_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0605_),
    .B(_0656_),
    .C(_0657_),
    .Y(_0658_)
);

sky130_fd_sc_hd__a21o_4 _1473_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0389_),
    .A2(_0590_),
    .B1(_0391_),
    .X(_0659_)
);

sky130_fd_sc_hd__o32ai_4 _1474_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0596_),
    .A2(_0654_),
    .A3(_0655_),
    .B1(_0658_),
    .B2(_0659_),
    .Y(_0035_)
);

sky130_fd_sc_hd__a2bb2o_4 _1475_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(\COUNT_BB_ZERO_MIN[7] ),
    .A2_N(_0403_),
    .B1(_0340_),
    .B2(_0406_),
    .X(_0660_)
);

sky130_fd_sc_hd__or2_4 _1476_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0355_),
    .B(_0397_),
    .X(_0661_)
);

sky130_fd_sc_hd__o21ai_4 _1477_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0347_),
    .A2(_0425_),
    .B1(_0661_),
    .Y(_0662_)
);

sky130_fd_sc_hd__or2_4 _1478_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0609_),
    .B(_0544_),
    .X(_0663_)
);

sky130_fd_sc_hd__o22a_4 _1479_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0304_),
    .A2(\COUNT_BB_ZERO[1] ),
    .B1(_0306_),
    .B2(\COUNT_BB_ZERO[0] ),
    .X(_0664_)
);

sky130_fd_sc_hd__and2_4 _1480_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0304_),
    .B(_0530_),
    .X(_0665_)
);

sky130_fd_sc_hd__o22a_4 _1481_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0500_),
    .A2(_0419_),
    .B1(_0664_),
    .B2(_0665_),
    .X(_0666_)
);

sky130_fd_sc_hd__a2bb2o_4 _1482_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0309_),
    .A2_N(_0412_),
    .B1(_0320_),
    .B2(_0536_),
    .X(_0667_)
);

sky130_fd_sc_hd__o22a_4 _1483_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0320_),
    .A2(_0536_),
    .B1(_0666_),
    .B2(_0667_),
    .X(_0668_)
);

sky130_fd_sc_hd__a21o_4 _1484_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0609_),
    .A2(_0544_),
    .B1(_0668_),
    .X(_0669_)
);

sky130_fd_sc_hd__a22oi_4 _1485_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0339_),
    .A2(_0400_),
    .B1(_0663_),
    .B2(_0669_),
    .Y(_0670_)
);

sky130_fd_sc_hd__a2111oi_4 _1486_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0347_),
    .A2(_0425_),
    .B1(_0660_),
    .C1(_0662_),
    .D1(_0670_),
    .Y(_0671_)
);

sky130_fd_sc_hd__a32o_4 _1487_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0399_),
    .A2(_0394_),
    .A3(_0661_),
    .B1(_0356_),
    .B2(_0397_),
    .X(_0672_)
);

sky130_fd_sc_hd__o22a_4 _1488_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0446_),
    .A2(_0428_),
    .B1(_0671_),
    .B2(_0672_),
    .X(_0673_)
);

sky130_fd_sc_hd__a2bb2o_4 _1489_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0364_),
    .A2_N(_0554_),
    .B1(_0373_),
    .B2(_0485_),
    .X(_0674_)
);

sky130_fd_sc_hd__o22a_4 _1490_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0374_),
    .A2(_0485_),
    .B1(_0673_),
    .B2(_0674_),
    .X(_0675_)
);

sky130_fd_sc_hd__a21o_4 _1491_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0387_),
    .A2(\COUNT_BB_ZERO[10] ),
    .B1(_0675_),
    .X(_0676_)
);

sky130_fd_sc_hd__o21a_4 _1492_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0388_),
    .A2(\COUNT_BB_ZERO[10] ),
    .B1(_0676_),
    .X(_0677_)
);

sky130_fd_sc_hd__o21a_4 _1493_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0415_),
    .A2(_0677_),
    .B1(_0069_),
    .X(_0023_)
);

sky130_fd_sc_hd__buf_1 _1494_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0145_),
    .X(_0678_)
);

sky130_fd_sc_hd__inv_8 _1495_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0677_),
    .Y(_0679_)
);

sky130_fd_sc_hd__buf_1 _1496_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0679_),
    .X(_0680_)
);

sky130_fd_sc_hd__or2_4 _1497_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0530_),
    .B(\COUNT_BB_ZERO[0] ),
    .X(_0681_)
);

sky130_fd_sc_hd__or2_4 _1498_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0413_),
    .B(_0415_),
    .X(_0682_)
);

sky130_fd_sc_hd__and4_4 _1499_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0678_),
    .B(_0680_),
    .C(_0681_),
    .D(_0682_),
    .X(_0025_)
);

sky130_fd_sc_hd__nand2_4 _1500_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0412_),
    .B(_0682_),
    .Y(_0683_)
);

sky130_fd_sc_hd__or2_4 _1501_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0412_),
    .B(_0682_),
    .X(_0684_)
);

sky130_fd_sc_hd__and4_4 _1502_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0678_),
    .B(_0680_),
    .C(_0683_),
    .D(_0684_),
    .X(_0026_)
);

sky130_fd_sc_hd__or2_4 _1503_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0411_),
    .B(_0684_),
    .X(_0685_)
);

sky130_fd_sc_hd__nand2_4 _1504_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0411_),
    .B(_0684_),
    .Y(_0686_)
);

sky130_fd_sc_hd__and4_4 _1505_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0678_),
    .B(_0680_),
    .C(_0685_),
    .D(_0686_),
    .X(_0027_)
);

sky130_fd_sc_hd__buf_1 _1506_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0307_),
    .X(_0687_)
);

sky130_fd_sc_hd__nand2_4 _1507_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0408_),
    .B(_0685_),
    .Y(_0688_)
);

sky130_fd_sc_hd__or2_4 _1508_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0408_),
    .B(_0685_),
    .X(_0689_)
);

sky130_fd_sc_hd__and4_4 _1509_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0687_),
    .B(_0680_),
    .C(_0688_),
    .D(_0689_),
    .X(_0028_)
);

sky130_fd_sc_hd__nand2_4 _1510_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0406_),
    .B(_0689_),
    .Y(_0690_)
);

sky130_fd_sc_hd__or2_4 _1511_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0406_),
    .B(_0689_),
    .X(_0691_)
);

sky130_fd_sc_hd__and4_4 _1512_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0687_),
    .B(_0680_),
    .C(_0690_),
    .D(_0691_),
    .X(_0029_)
);

sky130_fd_sc_hd__nand2_4 _1513_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0425_),
    .B(_0691_),
    .Y(_0692_)
);

sky130_fd_sc_hd__or2_4 _1514_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0425_),
    .B(_0691_),
    .X(_0693_)
);

sky130_fd_sc_hd__and4_4 _1515_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0687_),
    .B(_0679_),
    .C(_0692_),
    .D(_0693_),
    .X(_0030_)
);

sky130_fd_sc_hd__or2_4 _1516_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0403_),
    .B(_0693_),
    .X(_0694_)
);

sky130_fd_sc_hd__nand2_4 _1517_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0403_),
    .B(_0693_),
    .Y(_0695_)
);

sky130_fd_sc_hd__and4_4 _1518_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0687_),
    .B(_0679_),
    .C(_0694_),
    .D(_0695_),
    .X(_0031_)
);

sky130_fd_sc_hd__nand2_4 _1519_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0554_),
    .B(_0694_),
    .Y(_0696_)
);

sky130_fd_sc_hd__or2_4 _1520_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0554_),
    .B(_0694_),
    .X(_0697_)
);

sky130_fd_sc_hd__and4_4 _1521_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0687_),
    .B(_0679_),
    .C(_0696_),
    .D(_0697_),
    .X(_0032_)
);

sky130_fd_sc_hd__or2_4 _1522_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0528_),
    .B(_0697_),
    .X(_0698_)
);

sky130_fd_sc_hd__nand2_4 _1523_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0528_),
    .B(_0697_),
    .Y(_0699_)
);

sky130_fd_sc_hd__and4_4 _1524_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0307_),
    .B(_0679_),
    .C(_0698_),
    .D(_0699_),
    .X(_0033_)
);

sky130_fd_sc_hd__nor2_4 _1525_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0443_),
    .B(_0698_),
    .Y(_0700_)
);

sky130_fd_sc_hd__a2111oi_4 _1526_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0443_),
    .A2(_0698_),
    .B1(_0700_),
    .C1(_0272_),
    .D1(_0677_),
    .Y(_0024_)
);

sky130_fd_sc_hd__o21a_4 _1527_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0598_),
    .A2(_0677_),
    .B1(_0069_),
    .X(_0067_)
);

sky130_fd_sc_hd__inv_8 _1528_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ONE),
    .Y(_0701_)
);

sky130_fd_sc_hd__buf_1 _1529_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0701_),
    .X(_0702_)
);

sky130_fd_sc_hd__buf_1 _1530_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[9] ),
    .X(_0703_)
);

sky130_fd_sc_hd__buf_1 _1531_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0703_),
    .X(_0704_)
);

sky130_fd_sc_hd__buf_1 _1532_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[6] ),
    .X(_0705_)
);

sky130_fd_sc_hd__and2_4 _1533_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0360_),
    .B(_0705_),
    .X(_0706_)
);

sky130_fd_sc_hd__inv_8 _1534_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[8] ),
    .Y(_0707_)
);

sky130_fd_sc_hd__inv_8 _1535_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[6] ),
    .Y(_0708_)
);

sky130_fd_sc_hd__buf_1 _1536_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[5] ),
    .X(_0709_)
);

sky130_fd_sc_hd__a2bb2o_4 _1537_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0707_),
    .A2_N(\COUNT_BB_ONE[7] ),
    .B1(_0708_),
    .B2(_0709_),
    .X(_0710_)
);

sky130_fd_sc_hd__inv_8 _1538_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[7] ),
    .Y(_0711_)
);

sky130_fd_sc_hd__or2_4 _1539_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0368_),
    .B(_0711_),
    .X(_0712_)
);

sky130_fd_sc_hd__o21ai_4 _1540_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0360_),
    .A2(_0705_),
    .B1(_0712_),
    .Y(_0713_)
);

sky130_fd_sc_hd__inv_8 _1541_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[5] ),
    .Y(_0714_)
);

sky130_fd_sc_hd__inv_8 _1542_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[4] ),
    .Y(_0715_)
);

sky130_fd_sc_hd__or2_4 _1543_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0344_),
    .B(_0715_),
    .X(_0716_)
);

sky130_fd_sc_hd__inv_8 _1544_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[3] ),
    .Y(_0717_)
);

sky130_fd_sc_hd__inv_8 _1545_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[2] ),
    .Y(_0718_)
);

sky130_fd_sc_hd__inv_8 _1546_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[1] ),
    .Y(_0719_)
);

sky130_fd_sc_hd__inv_8 _1547_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[0] ),
    .Y(_0720_)
);

sky130_fd_sc_hd__buf_1 _1548_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0720_),
    .X(_0721_)
);

sky130_fd_sc_hd__o22a_4 _1549_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[2] ),
    .A2(_0719_),
    .B1(_0296_),
    .B2(_0721_),
    .X(_0722_)
);

sky130_fd_sc_hd__and2_4 _1550_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0314_),
    .B(_0719_),
    .X(_0723_)
);

sky130_fd_sc_hd__o22a_4 _1551_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0326_),
    .A2(_0718_),
    .B1(_0722_),
    .B2(_0723_),
    .X(_0724_)
);

sky130_fd_sc_hd__buf_1 _1552_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[2] ),
    .X(_0725_)
);

sky130_fd_sc_hd__a2bb2o_4 _1553_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0324_),
    .A2_N(_0725_),
    .B1(_0334_),
    .B2(_0717_),
    .X(_0726_)
);

sky130_fd_sc_hd__o22a_4 _1554_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0334_),
    .A2(_0717_),
    .B1(_0724_),
    .B2(_0726_),
    .X(_0727_)
);

sky130_fd_sc_hd__a21o_4 _1555_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0344_),
    .A2(_0715_),
    .B1(_0727_),
    .X(_0728_)
);

sky130_fd_sc_hd__a22oi_4 _1556_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[6] ),
    .A2(_0714_),
    .B1(_0716_),
    .B2(_0728_),
    .Y(_0729_)
);

sky130_fd_sc_hd__inv_8 _1557_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0705_),
    .Y(_0730_)
);

sky130_fd_sc_hd__buf_1 _1558_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0711_),
    .X(_0731_)
);

sky130_fd_sc_hd__a32oi_4 _1559_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[7] ),
    .A2(_0730_),
    .A3(_0712_),
    .B1(_0368_),
    .B2(_0731_),
    .Y(_0732_)
);

sky130_fd_sc_hd__o41a_4 _1560_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0706_),
    .A2(_0710_),
    .A3(_0713_),
    .A4(_0729_),
    .B1(_0732_),
    .X(_0733_)
);

sky130_fd_sc_hd__buf_1 _1561_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[8] ),
    .X(_0734_)
);

sky130_fd_sc_hd__a2bb2o_4 _1562_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0383_),
    .A2_N(_0703_),
    .B1(_0378_),
    .B2(_0734_),
    .X(_0735_)
);

sky130_fd_sc_hd__o22a_4 _1563_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0382_),
    .A2(_0703_),
    .B1(_0378_),
    .B2(_0734_),
    .X(_0736_)
);

sky130_fd_sc_hd__o21a_4 _1564_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0733_),
    .A2(_0735_),
    .B1(_0736_),
    .X(_0737_)
);

sky130_fd_sc_hd__a211o_4 _1565_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0383_),
    .A2(_0704_),
    .B1(\COUNT_BB_ONE[10] ),
    .C1(_0737_),
    .X(_0738_)
);

sky130_fd_sc_hd__inv_8 _1566_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0738_),
    .Y(_0739_)
);

sky130_fd_sc_hd__or4_4 _1567_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[8] ),
    .B(\COUNT_BB_ONE[7] ),
    .C(\COUNT_BB_ONE[6] ),
    .D(\COUNT_BB_ONE[5] ),
    .X(_0740_)
);

sky130_fd_sc_hd__or4_4 _1568_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[4] ),
    .B(\COUNT_BB_ONE[3] ),
    .C(\COUNT_BB_ONE[2] ),
    .D(\COUNT_BB_ONE[1] ),
    .X(_0741_)
);

sky130_fd_sc_hd__nor4_4 _1569_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[10] ),
    .B(\COUNT_BB_ONE[9] ),
    .C(_0740_),
    .D(_0741_),
    .Y(_0742_)
);

sky130_fd_sc_hd__and2_4 _1570_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0739_),
    .B(_0742_),
    .X(_0743_)
);

sky130_fd_sc_hd__or2_4 _1571_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0299_),
    .B(_0743_),
    .X(_0744_)
);

sky130_fd_sc_hd__buf_1 _1572_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0744_),
    .X(_0745_)
);

sky130_fd_sc_hd__inv_8 _1573_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0745_),
    .Y(_0746_)
);

sky130_fd_sc_hd__and2_4 _1574_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0299_),
    .B(_0743_),
    .X(_0747_)
);

sky130_fd_sc_hd__inv_8 _1575_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[10] ),
    .Y(_0748_)
);

sky130_fd_sc_hd__buf_1 _1576_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0748_),
    .X(_0749_)
);

sky130_fd_sc_hd__and2_4 _1577_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0377_),
    .B(_0444_),
    .X(_0750_)
);

sky130_fd_sc_hd__and2_4 _1578_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0707_),
    .B(_0447_),
    .X(_0751_)
);

sky130_fd_sc_hd__and2_4 _1579_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0359_),
    .B(_0449_),
    .X(_0752_)
);

sky130_fd_sc_hd__a2bb2o_4 _1580_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0708_),
    .A2_N(_0452_),
    .B1(_0708_),
    .B2(_0452_),
    .X(_0753_)
);

sky130_fd_sc_hd__or2_4 _1581_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[5] ),
    .B(SCAN_IN[5]),
    .X(_0754_)
);

sky130_fd_sc_hd__o21ai_4 _1582_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0343_),
    .A2(_0454_),
    .B1(_0754_),
    .Y(_0755_)
);

sky130_fd_sc_hd__inv_8 _1583_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[4] ),
    .Y(_0756_)
);

sky130_fd_sc_hd__a2bb2o_4 _1584_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0756_),
    .A2_N(_0459_),
    .B1(_0756_),
    .B2(_0459_),
    .X(_0757_)
);

sky130_fd_sc_hd__or2_4 _1585_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[3] ),
    .B(SCAN_IN[3]),
    .X(_0758_)
);

sky130_fd_sc_hd__o21ai_4 _1586_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0324_),
    .A2(_0461_),
    .B1(_0758_),
    .Y(_0759_)
);

sky130_fd_sc_hd__inv_8 _1587_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[2] ),
    .Y(_0760_)
);

sky130_fd_sc_hd__o22a_4 _1588_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0760_),
    .A2(_0465_),
    .B1(\COUNT_BB_ONE_MIN[2] ),
    .B2(SCAN_IN[2]),
    .X(_0761_)
);

sky130_fd_sc_hd__inv_8 _1589_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0761_),
    .Y(_0762_)
);

sky130_fd_sc_hd__o22a_4 _1590_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0298_),
    .A2(_0468_),
    .B1(\COUNT_BB_ONE_MIN[1] ),
    .B2(SCAN_IN[1]),
    .X(_0763_)
);

sky130_fd_sc_hd__and3_4 _1591_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[0] ),
    .B(SCAN_IN[0]),
    .C(_0763_),
    .X(_0764_)
);

sky130_fd_sc_hd__a21o_4 _1592_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[1] ),
    .A2(SCAN_IN[1]),
    .B1(_0764_),
    .X(_0765_)
);

sky130_fd_sc_hd__inv_8 _1593_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0765_),
    .Y(_0766_)
);

sky130_fd_sc_hd__nor3_4 _1594_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0759_),
    .B(_0762_),
    .C(_0766_),
    .Y(_0767_)
);

sky130_fd_sc_hd__a32o_4 _1595_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[2] ),
    .A2(SCAN_IN[2]),
    .A3(_0758_),
    .B1(\COUNT_BB_ONE_MIN[3] ),
    .B2(SCAN_IN[3]),
    .X(_0768_)
);

sky130_fd_sc_hd__nor2_4 _1596_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0767_),
    .B(_0768_),
    .Y(_0769_)
);

sky130_fd_sc_hd__nor3_4 _1597_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0755_),
    .B(_0757_),
    .C(_0769_),
    .Y(_0770_)
);

sky130_fd_sc_hd__a32o_4 _1598_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[4] ),
    .A2(SCAN_IN[4]),
    .A3(_0754_),
    .B1(\COUNT_BB_ONE_MIN[5] ),
    .B2(SCAN_IN[5]),
    .X(_0771_)
);

sky130_fd_sc_hd__nor2_4 _1599_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0770_),
    .B(_0771_),
    .Y(_0772_)
);

sky130_fd_sc_hd__o22a_4 _1600_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0708_),
    .A2(_0452_),
    .B1(_0753_),
    .B2(_0772_),
    .X(_0773_)
);

sky130_fd_sc_hd__o22a_4 _1601_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0360_),
    .A2(_0449_),
    .B1(_0752_),
    .B2(_0773_),
    .X(_0774_)
);

sky130_fd_sc_hd__o22a_4 _1602_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0707_),
    .A2(_0447_),
    .B1(_0751_),
    .B2(_0774_),
    .X(_0775_)
);

sky130_fd_sc_hd__o22a_4 _1603_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0378_),
    .A2(_0444_),
    .B1(_0750_),
    .B2(_0775_),
    .X(_0776_)
);

sky130_fd_sc_hd__o22a_4 _1604_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0383_),
    .A2(SCAN_IN[10]),
    .B1(\COUNT_BB_ONE_MIN[10] ),
    .B2(_0482_),
    .X(_0777_)
);

sky130_fd_sc_hd__xor2_4 _1605_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0776_),
    .B(_0777_),
    .X(_0778_)
);

sky130_fd_sc_hd__a21oi_4 _1606_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0368_),
    .A2(SCAN_IN[8]),
    .B1(_0751_),
    .Y(_0779_)
);

sky130_fd_sc_hd__xor2_4 _1607_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0774_),
    .B(_0779_),
    .X(_0780_)
);

sky130_fd_sc_hd__or2_4 _1608_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0734_),
    .B(_0780_),
    .X(_0781_)
);

sky130_fd_sc_hd__buf_1 _1609_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[7] ),
    .X(_0782_)
);

sky130_fd_sc_hd__a21o_4 _1610_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[7] ),
    .A2(SCAN_IN[7]),
    .B1(_0752_),
    .X(_0783_)
);

sky130_fd_sc_hd__a2bb2o_4 _1611_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0773_),
    .A2_N(_0783_),
    .B1(_0773_),
    .B2(_0783_),
    .X(_0784_)
);

sky130_fd_sc_hd__or2_4 _1612_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0782_),
    .B(_0784_),
    .X(_0785_)
);

sky130_fd_sc_hd__buf_1 _1613_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0717_),
    .X(_0786_)
);

sky130_fd_sc_hd__or2_4 _1614_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0766_),
    .B(_0762_),
    .X(_0787_)
);

sky130_fd_sc_hd__o21a_4 _1615_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0760_),
    .A2(_0465_),
    .B1(_0787_),
    .X(_0788_)
);

sky130_fd_sc_hd__a2bb2o_4 _1616_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0759_),
    .A2_N(_0788_),
    .B1(_0759_),
    .B2(_0788_),
    .X(_0789_)
);

sky130_fd_sc_hd__inv_8 _1617_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0789_),
    .Y(_0790_)
);

sky130_fd_sc_hd__inv_8 _1618_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0763_),
    .Y(_0791_)
);

sky130_fd_sc_hd__or2_4 _1619_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[0] ),
    .B(_0720_),
    .X(_0792_)
);

sky130_fd_sc_hd__and2_4 _1620_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[0] ),
    .B(_0720_),
    .X(_0793_)
);

sky130_fd_sc_hd__a21o_4 _1621_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[0]),
    .A2(_0792_),
    .B1(_0793_),
    .X(_0794_)
);

sky130_fd_sc_hd__a21oi_4 _1622_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0719_),
    .A2(_0763_),
    .B1(_0794_),
    .Y(_0795_)
);

sky130_fd_sc_hd__a211o_4 _1623_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE[1] ),
    .A2(_0791_),
    .B1(_0764_),
    .C1(_0795_),
    .X(_0796_)
);

sky130_fd_sc_hd__o21ai_4 _1624_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0765_),
    .A2(_0761_),
    .B1(_0787_),
    .Y(_0797_)
);

sky130_fd_sc_hd__a21oi_4 _1625_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0796_),
    .A2(_0797_),
    .B1(_0725_),
    .Y(_0798_)
);

sky130_fd_sc_hd__nor2_4 _1626_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0796_),
    .B(_0797_),
    .Y(_0799_)
);

sky130_fd_sc_hd__o22a_4 _1627_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0786_),
    .A2(_0790_),
    .B1(_0798_),
    .B2(_0799_),
    .X(_0800_)
);

sky130_fd_sc_hd__buf_1 _1628_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[3] ),
    .X(_0801_)
);

sky130_fd_sc_hd__a2bb2o_4 _1629_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0769_),
    .A2_N(_0757_),
    .B1(_0769_),
    .B2(_0757_),
    .X(_0802_)
);

sky130_fd_sc_hd__or2_4 _1630_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[4] ),
    .B(_0802_),
    .X(_0803_)
);

sky130_fd_sc_hd__o21ai_4 _1631_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0801_),
    .A2(_0789_),
    .B1(_0803_),
    .Y(_0804_)
);

sky130_fd_sc_hd__buf_1 _1632_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0756_),
    .X(_0805_)
);

sky130_fd_sc_hd__o22a_4 _1633_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0805_),
    .A2(_0459_),
    .B1(_0769_),
    .B2(_0757_),
    .X(_0806_)
);

sky130_fd_sc_hd__a2bb2o_4 _1634_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0755_),
    .A2_N(_0806_),
    .B1(_0755_),
    .B2(_0806_),
    .X(_0807_)
);

sky130_fd_sc_hd__buf_1 _1635_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[4] ),
    .X(_0808_)
);

sky130_fd_sc_hd__a22oi_4 _1636_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0709_),
    .A2(_0807_),
    .B1(_0808_),
    .B2(_0802_),
    .Y(_0809_)
);

sky130_fd_sc_hd__o21a_4 _1637_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0800_),
    .A2(_0804_),
    .B1(_0809_),
    .X(_0810_)
);

sky130_fd_sc_hd__buf_1 _1638_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0705_),
    .X(_0811_)
);

sky130_fd_sc_hd__a2bb2o_4 _1639_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0753_),
    .A2_N(_0772_),
    .B1(_0753_),
    .B2(_0772_),
    .X(_0812_)
);

sky130_fd_sc_hd__or2_4 _1640_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0709_),
    .B(_0807_),
    .X(_0813_)
);

sky130_fd_sc_hd__o21ai_4 _1641_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0811_),
    .A2(_0812_),
    .B1(_0813_),
    .Y(_0814_)
);

sky130_fd_sc_hd__a22oi_4 _1642_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0782_),
    .A2(_0784_),
    .B1(_0811_),
    .B2(_0812_),
    .Y(_0815_)
);

sky130_fd_sc_hd__o21ai_4 _1643_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0810_),
    .A2(_0814_),
    .B1(_0815_),
    .Y(_0816_)
);

sky130_fd_sc_hd__buf_1 _1644_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0734_),
    .X(_0817_)
);

sky130_fd_sc_hd__a32o_4 _1645_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0781_),
    .A2(_0785_),
    .A3(_0816_),
    .B1(_0817_),
    .B2(_0780_),
    .X(_0818_)
);

sky130_fd_sc_hd__nor2_4 _1646_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0704_),
    .B(_0818_),
    .Y(_0819_)
);

sky130_fd_sc_hd__a21o_4 _1647_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(\COUNT_BB_ONE_MIN[9] ),
    .A2(SCAN_IN[9]),
    .B1(_0750_),
    .X(_0820_)
);

sky130_fd_sc_hd__a2bb2oi_4 _1648_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0775_),
    .A2_N(_0820_),
    .B1(_0775_),
    .B2(_0820_),
    .Y(_0821_)
);

sky130_fd_sc_hd__a21boi_4 _1649_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0704_),
    .A2(_0818_),
    .B1_N(_0821_),
    .Y(_0822_)
);

sky130_fd_sc_hd__a211o_4 _1650_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0748_),
    .A2(_0778_),
    .B1(_0819_),
    .C1(_0822_),
    .X(_0823_)
);

sky130_fd_sc_hd__o21ai_4 _1651_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0749_),
    .A2(_0778_),
    .B1(_0823_),
    .Y(_0824_)
);

sky130_fd_sc_hd__inv_8 _1652_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0703_),
    .Y(_0825_)
);

sky130_fd_sc_hd__or2_4 _1653_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[20]),
    .B(_0825_),
    .X(_0826_)
);

sky130_fd_sc_hd__nor2_4 _1654_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[18]),
    .B(_0731_),
    .Y(_0827_)
);

sky130_fd_sc_hd__a2bb2o_4 _1655_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0547_),
    .A2_N(\COUNT_BB_ONE[6] ),
    .B1(SCAN_IN[18]),
    .B2(_0731_),
    .X(_0828_)
);

sky130_fd_sc_hd__a211o_4 _1656_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0547_),
    .A2(_0705_),
    .B1(_0827_),
    .C1(_0828_),
    .X(_0829_)
);

sky130_fd_sc_hd__and2_4 _1657_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[11]),
    .B(_0721_),
    .X(_0830_)
);

sky130_fd_sc_hd__buf_1 _1658_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0719_),
    .X(_0831_)
);

sky130_fd_sc_hd__and2_4 _1659_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[12]),
    .B(_0831_),
    .X(_0832_)
);

sky130_fd_sc_hd__and2_4 _1660_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[13]),
    .B(_0718_),
    .X(_0833_)
);

sky130_fd_sc_hd__a2111o_4 _1661_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0542_),
    .A2(\COUNT_BB_ONE[9] ),
    .B1(_0830_),
    .C1(_0832_),
    .D1(_0833_),
    .X(_0834_)
);

sky130_fd_sc_hd__or2_4 _1662_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[16]),
    .B(_0714_),
    .X(_0835_)
);

sky130_fd_sc_hd__buf_1 _1663_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0835_),
    .X(_0836_)
);

sky130_fd_sc_hd__inv_8 _1664_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0836_),
    .Y(_0837_)
);

sky130_fd_sc_hd__a2bb2o_4 _1665_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0560_),
    .A2_N(\COUNT_BB_ONE[5] ),
    .B1(SCAN_IN[15]),
    .B2(_0715_),
    .X(_0838_)
);

sky130_fd_sc_hd__a211o_4 _1666_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0543_),
    .A2(\COUNT_BB_ONE[4] ),
    .B1(_0837_),
    .C1(_0838_),
    .X(_0839_)
);

sky130_fd_sc_hd__o22a_4 _1667_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0558_),
    .A2(_0734_),
    .B1(_0542_),
    .B2(\COUNT_BB_ONE[9] ),
    .X(_0840_)
);

sky130_fd_sc_hd__inv_8 _1668_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[8] ),
    .Y(_0841_)
);

sky130_fd_sc_hd__or2_4 _1669_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SCAN_IN[14]),
    .B(_0786_),
    .X(_0842_)
);

sky130_fd_sc_hd__o21a_4 _1670_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[19]),
    .A2(_0841_),
    .B1(_0842_),
    .X(_0843_)
);

sky130_fd_sc_hd__o22a_4 _1671_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[12]),
    .A2(_0831_),
    .B1(SCAN_IN[11]),
    .B2(_0721_),
    .X(_0844_)
);

sky130_fd_sc_hd__o22a_4 _1672_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0537_),
    .A2(\COUNT_BB_ONE[3] ),
    .B1(SCAN_IN[13]),
    .B2(_0718_),
    .X(_0845_)
);

sky130_fd_sc_hd__nand4_4 _1673_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0840_),
    .B(_0843_),
    .C(_0844_),
    .D(_0845_),
    .Y(_0846_)
);

sky130_fd_sc_hd__or4_4 _1674_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0829_),
    .B(_0834_),
    .C(_0839_),
    .D(_0846_),
    .X(_0847_)
);

sky130_fd_sc_hd__and2_4 _1675_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0558_),
    .B(_0817_),
    .X(_0848_)
);

sky130_fd_sc_hd__inv_8 _1676_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0839_),
    .Y(_0849_)
);

sky130_fd_sc_hd__o21a_4 _1677_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0832_),
    .A2(_0844_),
    .B1(_0845_),
    .X(_0850_)
);

sky130_fd_sc_hd__a211o_4 _1678_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[14]),
    .A2(_0786_),
    .B1(_0833_),
    .C1(_0850_),
    .X(_0851_)
);

sky130_fd_sc_hd__a32oi_4 _1679_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0849_),
    .A2(_0842_),
    .A3(_0851_),
    .B1(_0836_),
    .B2(_0838_),
    .Y(_0852_)
);

sky130_fd_sc_hd__inv_8 _1680_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0828_),
    .Y(_0853_)
);

sky130_fd_sc_hd__o22a_4 _1681_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0829_),
    .A2(_0852_),
    .B1(_0853_),
    .B2(_0827_),
    .X(_0854_)
);

sky130_fd_sc_hd__o21ai_4 _1682_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0848_),
    .A2(_0854_),
    .B1(_0840_),
    .Y(_0855_)
);

sky130_fd_sc_hd__a32o_4 _1683_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0826_),
    .A2(_0847_),
    .A3(_0855_),
    .B1(SCAN_IN[21]),
    .B2(_0748_),
    .X(_0856_)
);

sky130_fd_sc_hd__o21a_4 _1684_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(SCAN_IN[21]),
    .A2(_0749_),
    .B1(_0856_),
    .X(_0857_)
);

sky130_fd_sc_hd__or2_4 _1685_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0824_),
    .B(_0857_),
    .X(_0858_)
);

sky130_fd_sc_hd__buf_1 _1686_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0858_),
    .X(_0859_)
);

sky130_fd_sc_hd__and2_4 _1687_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0299_),
    .B(_0859_),
    .X(_0860_)
);

sky130_fd_sc_hd__buf_1 _1688_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ONE),
    .X(_0861_)
);

sky130_fd_sc_hd__buf_1 _1689_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0857_),
    .X(_0862_)
);

sky130_fd_sc_hd__buf_1 _1690_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0824_),
    .X(_0863_)
);

sky130_fd_sc_hd__nor3_4 _1691_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[0] ),
    .B(_0862_),
    .C(_0863_),
    .Y(_0864_)
);

sky130_fd_sc_hd__or2_4 _1692_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0861_),
    .B(_0864_),
    .X(_0865_)
);

sky130_fd_sc_hd__o32ai_4 _1693_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0702_),
    .A2(_0746_),
    .A3(_0747_),
    .B1(_0860_),
    .B2(_0865_),
    .Y(_0012_)
);

sky130_fd_sc_hd__or3_4 _1694_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[1] ),
    .B(_0862_),
    .C(_0863_),
    .X(_0866_)
);

sky130_fd_sc_hd__nand2_4 _1695_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0298_),
    .B(_0859_),
    .Y(_0867_)
);

sky130_fd_sc_hd__buf_1 _1696_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0739_),
    .X(_0868_)
);

sky130_fd_sc_hd__o22a_4 _1697_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0296_),
    .A2(_0868_),
    .B1(_0298_),
    .B2(_0738_),
    .X(_0869_)
);

sky130_fd_sc_hd__nand2_4 _1698_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0745_),
    .B(_0869_),
    .Y(_0870_)
);

sky130_fd_sc_hd__o21a_4 _1699_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0745_),
    .A2(_0869_),
    .B1(_0861_),
    .X(_0871_)
);

sky130_fd_sc_hd__a32o_4 _1700_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0702_),
    .A2(_0866_),
    .A3(_0867_),
    .B1(_0870_),
    .B2(_0871_),
    .X(_0014_)
);

sky130_fd_sc_hd__and2_4 _1701_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0760_),
    .B(_0859_),
    .X(_0872_)
);

sky130_fd_sc_hd__nor3_4 _1702_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0725_),
    .B(_0862_),
    .C(_0863_),
    .Y(_0873_)
);

sky130_fd_sc_hd__or2_4 _1703_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0861_),
    .B(_0873_),
    .X(_0874_)
);

sky130_fd_sc_hd__buf_1 _1704_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0738_),
    .X(_0875_)
);

sky130_fd_sc_hd__or2_4 _1705_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0300_),
    .B(_0742_),
    .X(_0876_)
);

sky130_fd_sc_hd__or2_4 _1706_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0760_),
    .B(_0876_),
    .X(_0877_)
);

sky130_fd_sc_hd__inv_8 _1707_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0877_),
    .Y(_0878_)
);

sky130_fd_sc_hd__a21oi_4 _1708_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0760_),
    .A2(_0876_),
    .B1(_0878_),
    .Y(_0879_)
);

sky130_fd_sc_hd__or2_4 _1709_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0875_),
    .B(_0879_),
    .X(_0880_)
);

sky130_fd_sc_hd__buf_1 _1710_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(MULTIBIT_ONE),
    .X(_0881_)
);

sky130_fd_sc_hd__o21a_4 _1711_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0317_),
    .A2(_0868_),
    .B1(_0881_),
    .X(_0882_)
);

sky130_fd_sc_hd__a2bb2o_4 _1712_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0872_),
    .A2_N(_0874_),
    .B1(_0880_),
    .B2(_0882_),
    .X(_0015_)
);

sky130_fd_sc_hd__buf_1 _1713_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0861_),
    .X(_0883_)
);

sky130_fd_sc_hd__buf_1 _1714_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0857_),
    .X(_0884_)
);

sky130_fd_sc_hd__buf_1 _1715_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0824_),
    .X(_0885_)
);

sky130_fd_sc_hd__nor3_4 _1716_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0801_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0886_)
);

sky130_fd_sc_hd__and2_4 _1717_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0325_),
    .B(_0859_),
    .X(_0887_)
);

sky130_fd_sc_hd__or2_4 _1718_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0326_),
    .B(_0878_),
    .X(_0888_)
);

sky130_fd_sc_hd__or2_4 _1719_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0325_),
    .B(_0877_),
    .X(_0889_)
);

sky130_fd_sc_hd__buf_1 _1720_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0738_),
    .X(_0890_)
);

sky130_fd_sc_hd__a21oi_4 _1721_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0888_),
    .A2(_0889_),
    .B1(_0890_),
    .Y(_0891_)
);

sky130_fd_sc_hd__a21o_4 _1722_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0328_),
    .A2(_0890_),
    .B1(_0702_),
    .X(_0892_)
);

sky130_fd_sc_hd__o32ai_4 _1723_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0883_),
    .A2(_0886_),
    .A3(_0887_),
    .B1(_0891_),
    .B2(_0892_),
    .Y(_0016_)
);

sky130_fd_sc_hd__nor3_4 _1724_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0808_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0893_)
);

sky130_fd_sc_hd__buf_1 _1725_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0858_),
    .X(_0894_)
);

sky130_fd_sc_hd__and2_4 _1726_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0805_),
    .B(_0894_),
    .X(_0895_)
);

sky130_fd_sc_hd__buf_1 _1727_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0868_),
    .X(_0896_)
);

sky130_fd_sc_hd__nor2_4 _1728_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0337_),
    .B(_0896_),
    .Y(_0897_)
);

sky130_fd_sc_hd__or2_4 _1729_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0805_),
    .B(_0889_),
    .X(_0898_)
);

sky130_fd_sc_hd__inv_8 _1730_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0898_),
    .Y(_0899_)
);

sky130_fd_sc_hd__a21o_4 _1731_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0805_),
    .A2(_0889_),
    .B1(_0899_),
    .X(_0900_)
);

sky130_fd_sc_hd__a21o_4 _1732_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0896_),
    .A2(_0900_),
    .B1(_0702_),
    .X(_0901_)
);

sky130_fd_sc_hd__o32ai_4 _1733_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0883_),
    .A2(_0893_),
    .A3(_0895_),
    .B1(_0897_),
    .B2(_0901_),
    .Y(_0017_)
);

sky130_fd_sc_hd__nor3_4 _1734_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0709_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0902_)
);

sky130_fd_sc_hd__and2_4 _1735_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0343_),
    .B(_0894_),
    .X(_0903_)
);

sky130_fd_sc_hd__or2_4 _1736_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0344_),
    .B(_0899_),
    .X(_0904_)
);

sky130_fd_sc_hd__or2_4 _1737_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0343_),
    .B(_0898_),
    .X(_0905_)
);

sky130_fd_sc_hd__a21oi_4 _1738_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0904_),
    .A2(_0905_),
    .B1(_0890_),
    .Y(_0906_)
);

sky130_fd_sc_hd__a21o_4 _1739_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0346_),
    .A2(_0890_),
    .B1(_0702_),
    .X(_0907_)
);

sky130_fd_sc_hd__o32ai_4 _1740_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0883_),
    .A2(_0902_),
    .A3(_0903_),
    .B1(_0906_),
    .B2(_0907_),
    .Y(_0018_)
);

sky130_fd_sc_hd__buf_1 _1741_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0708_),
    .X(_0908_)
);

sky130_fd_sc_hd__and2_4 _1742_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0908_),
    .B(_0859_),
    .X(_0909_)
);

sky130_fd_sc_hd__nor3_4 _1743_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0811_),
    .B(_0862_),
    .C(_0863_),
    .Y(_0910_)
);

sky130_fd_sc_hd__or2_4 _1744_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0861_),
    .B(_0910_),
    .X(_0911_)
);

sky130_fd_sc_hd__or2_4 _1745_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0908_),
    .B(_0905_),
    .X(_0912_)
);

sky130_fd_sc_hd__a21boi_4 _1746_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0908_),
    .A2(_0905_),
    .B1_N(_0912_),
    .Y(_0913_)
);

sky130_fd_sc_hd__or2_4 _1747_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0875_),
    .B(_0913_),
    .X(_0914_)
);

sky130_fd_sc_hd__o21a_4 _1748_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0353_),
    .A2(_0868_),
    .B1(_0881_),
    .X(_0915_)
);

sky130_fd_sc_hd__a2bb2o_4 _1749_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0909_),
    .A2_N(_0911_),
    .B1(_0914_),
    .B2(_0915_),
    .X(_0019_)
);

sky130_fd_sc_hd__nor3_4 _1750_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0782_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0916_)
);

sky130_fd_sc_hd__and2_4 _1751_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0361_),
    .B(_0894_),
    .X(_0917_)
);

sky130_fd_sc_hd__and2_4 _1752_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0361_),
    .B(_0912_),
    .X(_0918_)
);

sky130_fd_sc_hd__or2_4 _1753_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0361_),
    .B(_0912_),
    .X(_0919_)
);

sky130_fd_sc_hd__buf_1 _1754_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0919_),
    .X(_0920_)
);

sky130_fd_sc_hd__inv_8 _1755_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0920_),
    .Y(_0921_)
);

sky130_fd_sc_hd__o21a_4 _1756_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0918_),
    .A2(_0921_),
    .B1(_0896_),
    .X(_0922_)
);

sky130_fd_sc_hd__a21o_4 _1757_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0363_),
    .A2(_0875_),
    .B1(_0701_),
    .X(_0070_)
);

sky130_fd_sc_hd__o32ai_4 _1758_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0883_),
    .A2(_0916_),
    .A3(_0917_),
    .B1(_0922_),
    .B2(_0070_),
    .Y(_0020_)
);

sky130_fd_sc_hd__nor3_4 _1759_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0817_),
    .B(_0862_),
    .C(_0863_),
    .Y(_0071_)
);

sky130_fd_sc_hd__buf_1 _1760_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0707_),
    .X(_0072_)
);

sky130_fd_sc_hd__and2_4 _1761_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0858_),
    .X(_0073_)
);

sky130_fd_sc_hd__nor3_4 _1762_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0881_),
    .B(_0071_),
    .C(_0073_),
    .Y(_0074_)
);

sky130_fd_sc_hd__or2_4 _1763_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0920_),
    .X(_0075_)
);

sky130_fd_sc_hd__inv_8 _1764_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0075_),
    .Y(_0076_)
);

sky130_fd_sc_hd__a21o_4 _1765_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0072_),
    .A2(_0920_),
    .B1(_0076_),
    .X(_0077_)
);

sky130_fd_sc_hd__o21a_4 _1766_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0371_),
    .A2(_0868_),
    .B1(MULTIBIT_ONE),
    .X(_0078_)
);

sky130_fd_sc_hd__a21boi_4 _1767_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0896_),
    .A2(_0077_),
    .B1_N(_0078_),
    .Y(_0079_)
);

sky130_fd_sc_hd__or2_4 _1768_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0074_),
    .B(_0079_),
    .X(_0021_)
);

sky130_fd_sc_hd__nor3_4 _1769_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0704_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0080_)
);

sky130_fd_sc_hd__and2_4 _1770_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0379_),
    .B(_0894_),
    .X(_0081_)
);

sky130_fd_sc_hd__and2_4 _1771_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0379_),
    .B(_0075_),
    .X(_0082_)
);

sky130_fd_sc_hd__and2_4 _1772_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE_MIN[9] ),
    .B(_0076_),
    .X(_0083_)
);

sky130_fd_sc_hd__o21a_4 _1773_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0082_),
    .A2(_0083_),
    .B1(_0896_),
    .X(_0084_)
);

sky130_fd_sc_hd__a21o_4 _1774_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0381_),
    .A2(_0875_),
    .B1(_0701_),
    .X(_0085_)
);

sky130_fd_sc_hd__o32ai_4 _1775_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0881_),
    .A2(_0080_),
    .A3(_0081_),
    .B1(_0084_),
    .B2(_0085_),
    .Y(_0022_)
);

sky130_fd_sc_hd__inv_8 _1776_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0856_),
    .Y(_0086_)
);

sky130_fd_sc_hd__and3_4 _1777_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0749_),
    .B(_0086_),
    .C(_0823_),
    .X(_0087_)
);

sky130_fd_sc_hd__and2_4 _1778_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0384_),
    .B(_0894_),
    .X(_0088_)
);

sky130_fd_sc_hd__and2_4 _1779_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0384_),
    .B(_0083_),
    .X(_0089_)
);

sky130_fd_sc_hd__nor2_4 _1780_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0384_),
    .B(_0083_),
    .Y(_0090_)
);

sky130_fd_sc_hd__nor3_4 _1781_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0890_),
    .B(_0089_),
    .C(_0090_),
    .Y(_0091_)
);

sky130_fd_sc_hd__a21o_4 _1782_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0385_),
    .A2(_0875_),
    .B1(_0701_),
    .X(_0092_)
);

sky130_fd_sc_hd__o32ai_4 _1783_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0881_),
    .A2(_0087_),
    .A3(_0088_),
    .B1(_0091_),
    .B2(_0092_),
    .Y(_0013_)
);

sky130_fd_sc_hd__o22a_4 _1784_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0072_),
    .A2(_0817_),
    .B1(_0379_),
    .B2(_0704_),
    .X(_0093_)
);

sky130_fd_sc_hd__and2_4 _1785_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0817_),
    .X(_0094_)
);

sky130_fd_sc_hd__nor2_4 _1786_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0793_),
    .B(_0094_),
    .Y(_0095_)
);

sky130_fd_sc_hd__o21a_4 _1787_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0296_),
    .A2(_0831_),
    .B1(_0792_),
    .X(_0096_)
);

sky130_fd_sc_hd__o22a_4 _1788_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0325_),
    .A2(_0801_),
    .B1(_0314_),
    .B2(_0718_),
    .X(_0097_)
);

sky130_fd_sc_hd__and4_4 _1789_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0093_),
    .B(_0095_),
    .C(_0096_),
    .D(_0097_),
    .X(_0098_)
);

sky130_fd_sc_hd__and2_4 _1790_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0361_),
    .B(_0782_),
    .X(_0099_)
);

sky130_fd_sc_hd__o22a_4 _1791_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0908_),
    .A2(_0811_),
    .B1(_0360_),
    .B2(_0782_),
    .X(_0100_)
);

sky130_fd_sc_hd__inv_8 _1792_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0100_),
    .Y(_0101_)
);

sky130_fd_sc_hd__a211o_4 _1793_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0908_),
    .A2(_0811_),
    .B1(_0099_),
    .C1(_0101_),
    .X(_0102_)
);

sky130_fd_sc_hd__and2_4 _1794_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0314_),
    .B(_0718_),
    .X(_0103_)
);

sky130_fd_sc_hd__and2_4 _1795_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0296_),
    .B(_0831_),
    .X(_0104_)
);

sky130_fd_sc_hd__and2_4 _1796_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0378_),
    .B(_0703_),
    .X(_0105_)
);

sky130_fd_sc_hd__a2111o_4 _1797_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0325_),
    .A2(_0801_),
    .B1(_0103_),
    .C1(_0104_),
    .D1(_0105_),
    .X(_0106_)
);

sky130_fd_sc_hd__or2_4 _1798_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0344_),
    .B(_0714_),
    .X(_0107_)
);

sky130_fd_sc_hd__buf_1 _1799_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0107_),
    .X(_0108_)
);

sky130_fd_sc_hd__inv_8 _1800_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0108_),
    .Y(_0109_)
);

sky130_fd_sc_hd__a2bb2o_4 _1801_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0343_),
    .A2_N(_0709_),
    .B1(_0334_),
    .B2(_0715_),
    .X(_0110_)
);

sky130_fd_sc_hd__a211o_4 _1802_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0805_),
    .A2(_0808_),
    .B1(_0109_),
    .C1(_0110_),
    .X(_0111_)
);

sky130_fd_sc_hd__nor3_4 _1803_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0102_),
    .B(_0106_),
    .C(_0111_),
    .Y(_0112_)
);

sky130_fd_sc_hd__inv_8 _1804_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0111_),
    .Y(_0113_)
);

sky130_fd_sc_hd__or2_4 _1805_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0326_),
    .B(_0786_),
    .X(_0114_)
);

sky130_fd_sc_hd__o21a_4 _1806_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0104_),
    .A2(_0096_),
    .B1(_0097_),
    .X(_0115_)
);

sky130_fd_sc_hd__a211o_4 _1807_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0326_),
    .A2(_0786_),
    .B1(_0103_),
    .C1(_0115_),
    .X(_0116_)
);

sky130_fd_sc_hd__a32oi_4 _1808_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0113_),
    .A2(_0114_),
    .A3(_0116_),
    .B1(_0108_),
    .B2(_0110_),
    .Y(_0117_)
);

sky130_fd_sc_hd__o22a_4 _1809_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0102_),
    .A2(_0117_),
    .B1(_0100_),
    .B2(_0099_),
    .X(_0118_)
);

sky130_fd_sc_hd__o21a_4 _1810_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0094_),
    .A2(_0118_),
    .B1(_0093_),
    .X(_0119_)
);

sky130_fd_sc_hd__a211o_4 _1811_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0098_),
    .A2(_0112_),
    .B1(_0105_),
    .C1(_0119_),
    .X(_0120_)
);

sky130_fd_sc_hd__nor2_4 _1812_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0383_),
    .B(_0120_),
    .Y(_0121_)
);

sky130_fd_sc_hd__a2bb2o_4 _1813_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1_N(_0749_),
    .A2_N(_0121_),
    .B1(_0384_),
    .B2(_0120_),
    .X(_0122_)
);

sky130_fd_sc_hd__o21a_4 _1814_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0721_),
    .A2(_0122_),
    .B1(_0323_),
    .X(_0001_)
);

sky130_fd_sc_hd__and2_4 _1815_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[1] ),
    .B(\COUNT_BB_ONE[0] ),
    .X(_0123_)
);

sky130_fd_sc_hd__buf_1 _1816_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .X(_0124_)
);

sky130_fd_sc_hd__a2111oi_4 _1817_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0831_),
    .A2(_0721_),
    .B1(_0313_),
    .C1(_0123_),
    .D1(_0124_),
    .Y(_0003_)
);

sky130_fd_sc_hd__and2_4 _1818_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0725_),
    .B(_0123_),
    .X(_0125_)
);

sky130_fd_sc_hd__nor2_4 _1819_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0725_),
    .B(_0123_),
    .Y(_0126_)
);

sky130_fd_sc_hd__nor4_4 _1820_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0338_),
    .B(_0125_),
    .C(_0126_),
    .D(_0124_),
    .Y(_0004_)
);

sky130_fd_sc_hd__nor2_4 _1821_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0801_),
    .B(_0125_),
    .Y(_0127_)
);

sky130_fd_sc_hd__and2_4 _1822_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[3] ),
    .B(_0125_),
    .X(_0128_)
);

sky130_fd_sc_hd__nor4_4 _1823_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0338_),
    .B(_0127_),
    .C(_0128_),
    .D(_0124_),
    .Y(_0005_)
);

sky130_fd_sc_hd__nand2_4 _1824_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0808_),
    .B(_0128_),
    .Y(_0129_)
);

sky130_fd_sc_hd__or2_4 _1825_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0808_),
    .B(_0128_),
    .X(_0130_)
);

sky130_fd_sc_hd__inv_8 _1826_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .Y(_0131_)
);

sky130_fd_sc_hd__and4_4 _1827_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0329_),
    .B(_0129_),
    .C(_0130_),
    .D(_0131_),
    .X(_0006_)
);

sky130_fd_sc_hd__or2_4 _1828_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0714_),
    .B(_0129_),
    .X(_0132_)
);

sky130_fd_sc_hd__nand2_4 _1829_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0714_),
    .B(_0129_),
    .Y(_0133_)
);

sky130_fd_sc_hd__and4_4 _1830_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0329_),
    .B(_0132_),
    .C(_0133_),
    .D(_0131_),
    .X(_0007_)
);

sky130_fd_sc_hd__or2_4 _1831_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0730_),
    .B(_0132_),
    .X(_0134_)
);

sky130_fd_sc_hd__nand2_4 _1832_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0730_),
    .B(_0132_),
    .Y(_0135_)
);

sky130_fd_sc_hd__and4_4 _1833_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0294_),
    .B(_0134_),
    .C(_0135_),
    .D(_0131_),
    .X(_0008_)
);

sky130_fd_sc_hd__nand2_4 _1834_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0731_),
    .B(_0134_),
    .Y(_0136_)
);

sky130_fd_sc_hd__or2_4 _1835_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0731_),
    .B(_0134_),
    .X(_0137_)
);

sky130_fd_sc_hd__and4_4 _1836_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0294_),
    .B(_0136_),
    .C(_0137_),
    .D(_0131_),
    .X(_0009_)
);

sky130_fd_sc_hd__or2_4 _1837_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0841_),
    .B(_0137_),
    .X(_0138_)
);

sky130_fd_sc_hd__nand2_4 _1838_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0841_),
    .B(_0137_),
    .Y(_0139_)
);

sky130_fd_sc_hd__and4_4 _1839_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0294_),
    .B(_0138_),
    .C(_0139_),
    .D(_0131_),
    .X(_0010_)
);

sky130_fd_sc_hd__or2_4 _1840_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0825_),
    .B(_0138_),
    .X(_0140_)
);

sky130_fd_sc_hd__buf_1 _1841_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0140_),
    .X(_0141_)
);

sky130_fd_sc_hd__inv_8 _1842_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0141_),
    .Y(_0142_)
);

sky130_fd_sc_hd__a2111oi_4 _1843_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0825_),
    .A2(_0138_),
    .B1(_0678_),
    .C1(_0142_),
    .D1(_0124_),
    .Y(_0011_)
);

sky130_fd_sc_hd__and2_4 _1844_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(\COUNT_BB_ONE[10] ),
    .B(_0142_),
    .X(_0143_)
);

sky130_fd_sc_hd__a2111oi_4 _1845_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0749_),
    .A2(_0141_),
    .B1(_0678_),
    .C1(_0143_),
    .D1(_0124_),
    .Y(_0002_)
);

sky130_fd_sc_hd__inv_8 _1846_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(BB_IN),
    .Y(_0068_)
);

sky130_fd_sc_hd__or2_4 _1847_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(RESET_LIFTED_N),
    .B(RESET_LIFTED_P),
    .X(RESET_LIFTED)
);

sky130_fd_sc_hd__o21a_4 _1848_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0883_),
    .A2(_0122_),
    .B1(_0272_),
    .X(_0066_)
);

sky130_fd_sc_hd__conb_1 _1849_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .HI(_0923_)
);

sky130_fd_sc_hd__conb_1 _1850_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .HI(_0924_)
);

sky130_fd_sc_hd__dfrtp_4 _1851_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0000_),
    .Q(CLK_OUT),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1852_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0055_),
    .Q(\DIVISOR_COUNT[0] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1853_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0057_),
    .Q(\DIVISOR_COUNT[1] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1854_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0058_),
    .Q(\DIVISOR_COUNT[2] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1855_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0059_),
    .Q(\DIVISOR_COUNT[3] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1856_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0060_),
    .Q(\DIVISOR_COUNT[4] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1857_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0061_),
    .Q(\DIVISOR_COUNT[5] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1858_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0062_),
    .Q(\DIVISOR_COUNT[6] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1859_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0063_),
    .Q(\DIVISOR_COUNT[7] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1860_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0064_),
    .Q(\DIVISOR_COUNT[8] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1861_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0065_),
    .Q(\DIVISOR_COUNT[9] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1862_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0056_),
    .Q(\DIVISOR_COUNT[10] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1863_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0069_),
    .Q(ONE_CHECKED),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfrtp_4 _1864_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(P_CLK),
    .Q(ZERO_CHECKED),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfstp_4 _1865_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0046_),
    .Q(\COUNT_MIN[0] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfstp_4 _1866_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0047_),
    .Q(\COUNT_MIN[1] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__dfstp_4 _1867_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0048_),
    .Q(\COUNT_MIN[2] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1868_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0049_),
    .Q(\COUNT_MIN[3] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1869_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0050_),
    .Q(\COUNT_MIN[4] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1870_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0051_),
    .Q(\COUNT_MIN[5] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1871_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0052_),
    .Q(\COUNT_MIN[6] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1872_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0053_),
    .Q(\COUNT_MIN[7] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1873_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0054_),
    .Q(\COUNT_MIN[8] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfstp_4 _1874_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0045_),
    .Q(\COUNT_MIN[9] ),
    .SET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1875_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0034_),
    .Q(\COUNT_BB_ZERO_MIN[0] ),
    .RESET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1876_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0036_),
    .Q(\COUNT_BB_ZERO_MIN[1] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1877_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0037_),
    .Q(\COUNT_BB_ZERO_MIN[2] ),
    .RESET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1878_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0038_),
    .Q(\COUNT_BB_ZERO_MIN[3] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1879_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0039_),
    .Q(\COUNT_BB_ZERO_MIN[4] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1880_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0040_),
    .Q(\COUNT_BB_ZERO_MIN[5] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1881_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0041_),
    .Q(\COUNT_BB_ZERO_MIN[6] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1882_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0042_),
    .Q(\COUNT_BB_ZERO_MIN[7] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1883_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0043_),
    .Q(\COUNT_BB_ZERO_MIN[8] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1884_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0044_),
    .Q(\COUNT_BB_ZERO_MIN[9] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1885_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0035_),
    .Q(\COUNT_BB_ZERO_MIN[10] ),
    .SET_B(RESET_LIFTED),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1886_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0023_),
    .Q(\COUNT_BB_ZERO[0] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1887_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0025_),
    .Q(\COUNT_BB_ZERO[1] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1888_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0026_),
    .Q(\COUNT_BB_ZERO[2] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1889_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0027_),
    .Q(\COUNT_BB_ZERO[3] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1890_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0028_),
    .Q(\COUNT_BB_ZERO[4] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1891_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0029_),
    .Q(\COUNT_BB_ZERO[5] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1892_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0030_),
    .Q(\COUNT_BB_ZERO[6] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1893_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0031_),
    .Q(\COUNT_BB_ZERO[7] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__dfrtp_4 _1894_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0032_),
    .Q(\COUNT_BB_ZERO[8] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1895_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0033_),
    .Q(\COUNT_BB_ZERO[9] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1896_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0024_),
    .Q(\COUNT_BB_ZERO[10] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1897_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0067_),
    .Q(MULTIBIT_ZERO),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1898_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0012_),
    .Q(\COUNT_BB_ONE_MIN[0] ),
    .RESET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1899_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0014_),
    .Q(\COUNT_BB_ONE_MIN[1] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1900_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0015_),
    .Q(\COUNT_BB_ONE_MIN[2] ),
    .RESET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1901_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0016_),
    .Q(\COUNT_BB_ONE_MIN[3] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1902_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0017_),
    .Q(\COUNT_BB_ONE_MIN[4] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1903_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0018_),
    .Q(\COUNT_BB_ONE_MIN[5] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1904_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0019_),
    .Q(\COUNT_BB_ONE_MIN[6] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1905_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0020_),
    .Q(\COUNT_BB_ONE_MIN[7] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1906_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0021_),
    .Q(\COUNT_BB_ONE_MIN[8] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1907_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0022_),
    .Q(\COUNT_BB_ONE_MIN[9] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfstp_4 _1908_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0013_),
    .Q(\COUNT_BB_ONE_MIN[10] ),
    .SET_B(RESET_LIFTED),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1909_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0001_),
    .Q(\COUNT_BB_ONE[0] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1910_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0003_),
    .Q(\COUNT_BB_ONE[1] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1911_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0004_),
    .Q(\COUNT_BB_ONE[2] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1912_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0005_),
    .Q(\COUNT_BB_ONE[3] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1913_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0006_),
    .Q(\COUNT_BB_ONE[4] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1914_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0007_),
    .Q(\COUNT_BB_ONE[5] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1915_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0008_),
    .Q(\COUNT_BB_ONE[6] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1916_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0009_),
    .Q(\COUNT_BB_ONE[7] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1917_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0010_),
    .Q(\COUNT_BB_ONE[8] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1918_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0011_),
    .Q(\COUNT_BB_ONE[9] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1919_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0002_),
    .Q(\COUNT_BB_ONE[10] ),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1920_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0066_),
    .Q(MULTIBIT_ONE),
    .RESET_B(RESET_LIFTED),
    .CLK(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__dfrtp_4 _1921_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0923_),
    .Q(RESET_LIFTED_N),
    .RESET_B(RESET_N),
    .CLK(N_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1922_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0924_),
    .Q(RESET_LIFTED_P),
    .RESET_B(RESET_N),
    .CLK(P_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1923_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(BB_IN),
    .Q(P_CLK),
    .RESET_B(RESET_N),
    .CLK(clknet_1_0_0_clk_0_48)
);

sky130_fd_sc_hd__dfrtp_4 _1924_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0068_),
    .Q(N_CLK),
    .RESET_B(RESET_N),
    .CLK(clknet_1_1_0_clk_0_48)
);

sky130_fd_sc_hd__dfrtp_4 _1925_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(BB_IN),
    .Q(DATA_OUT),
    .RESET_B(RESET_N),
    .CLK(CLK_OUT)
);

sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_1_0_0_clk_1_0),
    .X(clk_0_0)
);

sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_16 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_1_1_0_clk_1_0),
    .X(clk_0_16)
);

sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_32 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_1_1_0_clk_1_0),
    .X(clk_0_32)
);

sky130_fd_sc_hd__clkbuf_4 _CTS_buf_1_48 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_1_0_0_clk_1_0),
    .X(clk_0_48)
);

sky130_fd_sc_hd__clkbuf_16 _CTS_root (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(CLK_IN),
    .X(clk_1_0)
);

sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_96 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_0_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clk_0_0),
    .X(clknet_0_clk_0_0)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk_0_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_0),
    .X(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk_0_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_0),
    .X(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_0_16 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clk_0_16),
    .X(clknet_0_clk_0_16)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_0_16 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_16),
    .X(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk_0_16 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_16),
    .X(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_0_32 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clk_0_32),
    .X(clknet_0_clk_0_32)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_0_32 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_32),
    .X(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk_0_32 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_32),
    .X(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_0_48 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clk_0_48),
    .X(clknet_0_clk_0_48)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk_0_48 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_48),
    .X(clknet_1_0_0_clk_0_48)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk_0_48 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_0_48),
    .X(clknet_1_1_0_clk_0_48)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_1_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clk_1_0),
    .X(clknet_0_clk_1_0)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk_1_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_1_0),
    .X(clknet_1_0_0_clk_1_0)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk_1_0 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_clk_1_0),
    .X(clknet_1_1_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1925__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(BB_IN)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1923__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(BB_IN)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1846__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(BB_IN)
);

sky130_fd_sc_hd__diode_2 ANTENNA__CTS_root_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK_IN)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1925__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK_OUT)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1087__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK_OUT)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1083__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK_OUT)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1066__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK_OUT)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1925__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1924__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1923__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1922__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1921__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1621__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1591__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1311__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1271__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1604__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1287__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1286__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1671__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1657__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1350__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1337__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1671__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1659__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1336__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1335__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1672__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1660__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1339__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1678__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1341__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1665__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1347__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1662__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1364__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1361__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1351__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1655__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1654__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1355__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1352__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1670__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1362__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1359__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1592__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1590__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1275__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1273__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1272__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1653__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1346__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1333__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1684__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1683__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1376__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1375__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1595__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1588__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1277__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1269__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1595__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1585__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1277__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1266__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1265__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1598__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1280__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1262__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1598__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1581__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1280__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1259__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1258__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1255__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1610__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1292__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1253__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1606__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1290__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1251__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1647__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1327__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1248__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SCAN_IN[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1815__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1691__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1547__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1844__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1575__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1569__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1565__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1815__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1623__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1568__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1546__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1568__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1552__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1545__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1822__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1672__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1628__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1568__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1544__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1666__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1635__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1630__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1568__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1542__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1665__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1567__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1541__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1536__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1655__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1567__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1532__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1609__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1567__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1538__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1537__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1668__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1567__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1561__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1667__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1661__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1569__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1530__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1620__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1619__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1591__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1092__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1090__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1604__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1188__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1185__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1592__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1590__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1091__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1089__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1595__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1588__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1587__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1549__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1108__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1595__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1585__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1122__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1598__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1583__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1131__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1598__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1581__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1142__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1141__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1556__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1535__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1152__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1559__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1162__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1159__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1169__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1772__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1647__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1182__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1179__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ONE_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1497__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1479__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1383__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1218__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1492__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1491__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1246__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1240__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1236__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1479__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1334__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1314__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1239__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1217__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1315__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1239__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1223__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1216__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1340__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1239__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1214__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1348__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1239__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1211__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1301__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1300__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1238__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1204__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1355__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1238__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1228__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1198__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1294__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1238__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1206__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1201__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1363__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1358__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1323__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1238__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1232__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1363__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1357__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1240__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1197__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1311__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1271__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1098__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1095__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1287__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1192__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1189__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1096__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1094__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1277__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1268__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1103__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1266__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1114__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1261__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1127__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1280__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1259__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1138__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1137__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1202__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1146__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1475__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1292__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1230__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1157__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1154__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1290__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1200__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1165__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1463__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1327__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1177__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1174__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_BB_ZERO_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0959__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1080__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0960__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1078__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1074__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0958__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1073__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1073__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0930__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1078__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1067__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0945__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0931__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1070__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1068__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1074__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1071__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0933__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1072__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1069__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0934__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1076__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1072__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0935__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1079__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0937__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0928__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\COUNT_MIN[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1080__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0964__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[0] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[10] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0965__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[1] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1019__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[2] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1023__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0955__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[3] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0943__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[4] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1033__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0946__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[5] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[6] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1077__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0973__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[7] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1079__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0988__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[8] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1077__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1053__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__0939__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(\DIVISOR_COUNT[9] )
);

sky130_fd_sc_hd__diode_2 ANTENNA__1766__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ONE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1710__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ONE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ONE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ONE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1457__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ZERO)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1402__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ZERO)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1380__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ZERO)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1195__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(MULTIBIT_ZERO)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1921__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1908__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1907__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1906__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1905__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1904__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1903__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1902__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1901__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1900__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1899__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1898__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(N_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0925__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(ONE_CHECKED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1922__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1885__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1884__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1883__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1882__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1881__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1880__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1879__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1878__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1877__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1876__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1875__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1864__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1126__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1119__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1086__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1064__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(P_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1920__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1919__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1918__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1917__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1916__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1915__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1914__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1913__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1912__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1911__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1910__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1909__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1908__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1907__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1906__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1905__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1904__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1903__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1902__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1901__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1900__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1899__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1898__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1897__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1896__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1895__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1894__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1893__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1892__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1891__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1890__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1889__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1888__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1887__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1886__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1885__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1884__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1883__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1882__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1881__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1880__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1879__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1878__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1877__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1876__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1875__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1874__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1873__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1872__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1871__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1870__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1869__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1868__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1867__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1866__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1865__SET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1864__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1863__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1862__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1861__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1860__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1859__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1858__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1857__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1856__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1855__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1854__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1853__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1852__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1851__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1847__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED_N)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1847__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET_LIFTED_P)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1065__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(ZERO_CHECKED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(ZERO_CHECKED)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1851__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0000_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1909__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0001_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1919__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0002_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1910__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0003_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1911__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0004_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1912__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0005_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1913__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0006_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1914__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0007_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1915__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0008_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1916__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0009_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1917__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0010_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1918__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0011_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1898__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0012_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1908__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1899__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0014_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1900__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1901__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1902__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1903__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0018_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1904__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1905__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0020_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1906__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0021_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1907__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0022_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1886__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0023_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1896__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0024_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1887__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0025_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1888__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0026_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1889__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0027_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1890__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1891__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0029_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1892__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0030_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1893__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1894__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1895__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0033_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1875__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1885__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0035_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1876__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0036_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1877__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0037_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1878__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0038_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1879__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1880__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1881__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0041_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1882__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0042_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1883__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1884__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0044_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1874__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1865__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1866__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0047_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1867__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0048_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1868__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1869__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0050_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1870__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0051_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1871__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0052_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1872__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1873__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1852__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0055_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1862__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0056_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1853__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0057_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1854__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0058_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1855__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1856__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0060_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1857__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0061_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1858__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0062_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1859__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0063_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1860__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1861__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0065_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1920__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0066_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1897__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0067_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1924__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1863__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1527__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1493__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1194__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1125__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1758__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0070_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1762__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0071_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1784__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1765__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1763__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1761__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1762__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0073_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0074_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1771__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0075_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1764__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0075_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1772__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0076_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1765__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0076_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1767__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1767__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0078_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1768__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0079_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1775__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0080_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1775__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1773__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1780__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1779__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1773__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1775__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1775__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1777__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0086_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1783__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0087_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1783__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1781__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1781__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1783__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0091_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1783__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1810__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1789__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1810__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0094_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1786__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0094_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1789__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0095_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1806__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1789__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1806__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1789__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1811__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1809__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1793__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1809__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1792__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1793__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1809__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1803__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1807__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0103_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1797__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0103_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1806__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0104_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1797__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0104_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1811__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1797__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1803__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1799__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1808__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1800__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1802__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1808__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0110_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1802__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0110_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1804__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1803__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1811__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1808__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1808__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0114_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1807__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1808__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1809__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0117_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1810__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0118_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1811__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0119_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1813__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0120_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1812__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0120_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1813__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1848__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1826__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1816__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1814__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1819__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1818__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1817__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1845__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1843__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1823__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1820__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1817__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1822__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0125_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1821__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0125_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1820__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0125_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1820__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1823__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1825__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1824__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1823__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1829__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1828__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1827__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1827__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1839__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1836__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1833__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1830__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1827__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1832__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0132_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1831__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0132_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1830__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0132_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1830__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0133_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1835__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0134_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1834__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0134_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1833__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0134_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1833__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1836__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1838__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0137_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1837__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0137_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1836__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0137_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1843__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1840__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1839__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1839__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1841__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1845__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0141_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0141_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1844__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0142_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1843__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0142_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1845__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0143_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1087__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0144_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1085__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0144_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0144_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1494__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1107__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1100__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1063__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0146_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0146_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1079__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0147_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0147_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0148_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0148_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0930__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0148_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0945__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0931__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0945__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0151_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0151_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0933__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0151_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0152_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0152_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0934__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0152_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0153_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0153_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0935__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0153_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0937__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0936__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0156_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0156_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0983__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0156_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0156_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0940__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0157_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0939__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0157_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0158_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0158_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0941__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0159_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0942__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0161_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0951__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0944__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1070__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1068__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1031__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1027__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0164_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0951__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0164_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0950__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0165_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0948__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0165_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0166_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0948__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0166_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0949__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0167_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1005__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0168_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0168_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1074__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1071__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1038__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1034__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1004__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0173_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0955__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0173_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0956__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0174_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0175_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0957__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0175_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0176_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0177_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0178_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0961__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0178_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1080__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0179_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0961__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0179_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0180_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0180_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0181_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0181_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0999__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0183_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0183_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0968__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0967__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0968__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0967__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0186_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0187_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0188_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0188_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0189_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0190_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0972__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0190_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0191_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0981__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0192_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0192_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1072__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1048__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1046__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1045__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0981__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0194_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0976__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0194_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0195_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0195_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0196_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1040__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0980__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0200_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0200_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1001__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0201_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0201_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0984__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0202_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0203_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0203_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0204_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0205_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1077__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1062__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1061__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0992__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0207_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0989__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0207_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1079__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1054__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1052__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1051__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0991__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0992__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0209_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0209_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0210_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0210_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0993__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0211_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1000__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0212_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0212_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0213_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1082__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0214_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1037__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0214_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0214_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0997__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1032__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0216_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1030__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0216_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0998__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0216_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1080__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1011__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0219_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0220_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0221_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0222_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0227_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0228_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1035__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1012__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1011__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1017__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0230_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0230_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1037__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0231_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1030__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0231_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0231_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0232_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1078__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1074__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1021__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0234_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0234_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0235_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1073__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1073__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1025__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0237_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1024__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0237_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0237_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0238_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1078__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1067__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1027__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1025__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1031__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0242_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1034__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0243_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1029__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0243_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1033__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0244_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1030__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0244_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1031__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0245_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1059__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1051__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1049__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1042__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1039__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1036__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0247_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1044__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0248_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1041__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0248_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1036__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0248_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1057__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1050__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1041__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1036__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1039__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0250_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1060__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0251_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1058__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0251_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1048__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0251_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1038__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0251_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1039__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0252_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1072__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1069__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1044__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1043__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1042__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1043__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0254_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1042__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0254_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1043__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0255_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1046__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0256_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1045__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0256_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1054__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0257_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1050__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0257_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1046__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0257_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1047__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0258_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0259_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1049__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0260_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1052__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0261_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1051__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0261_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1052__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0262_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1060__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0263_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1058__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0263_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1056__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0263_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1055__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0264_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1060__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0265_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1056__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0265_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1057__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0266_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1059__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0267_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1059__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0268_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1062__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0269_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1061__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0269_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1063__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0270_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1063__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0271_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1848__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1526__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1112__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1102__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1088__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1084__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0273_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1066__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0273_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1088__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0274_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1069__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0275_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1069__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0276_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1082__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0277_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1071__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0278_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1075__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0279_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1075__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0280_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1075__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0281_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1075__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1082__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0283_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1077__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0284_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1081__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1081__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0286_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1081__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0287_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1081__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0288_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1082__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0289_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1083__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0290_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1085__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1084__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1088__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0292_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1088__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1836__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1833__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1193__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1087__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1088__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0295_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1795__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1787__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1697__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1549__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1090__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1111__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0297_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1109__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0297_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1102__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0297_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1697__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0298_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1695__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0298_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1590__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0298_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1093__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0298_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0299_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1574__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0299_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1571__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0299_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1093__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0299_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1705__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0300_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1102__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0300_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1389__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1275__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1273__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1220__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1095__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1106__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0302_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1104__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0302_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1102__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0302_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1397__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0303_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1273__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0303_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0303_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1480__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1479__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1389__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1387__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1101__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1397__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0305_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1099__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0305_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1479__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1379__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1245__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1242__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1101__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1524__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1506__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1136__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1113__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1101__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1102__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0308_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1482__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1221__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1220__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1106__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1104__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1117__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0310_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1105__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0310_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1118__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0311_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1106__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0311_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1403__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0312_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1112__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0312_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1817__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1173__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1153__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1135__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1112__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1794__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1788__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1550__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1111__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1109__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1123__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0315_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1110__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0315_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1124__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0316_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1111__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0316_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1711__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0317_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1112__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0317_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1410__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1277__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1222__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1117__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1115__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1267__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0319_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1224__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0319_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1116__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0319_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1483__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1482__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1411__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1118__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1130__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0321_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1128__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0321_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1118__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0321_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1414__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0322_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1125__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0322_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1814__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1184__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1164__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1145__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1125__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1586__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0324_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1553__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0324_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1121__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0324_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1797__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1788__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1719__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1717__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1124__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1807__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1805__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1718__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1551__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1123__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1134__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0327_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1132__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0327_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1124__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0327_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1722__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0328_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1125__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0328_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1830__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1827__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1173__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1153__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1135__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1280__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1225__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1224__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1130__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1128__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1139__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0331_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1129__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0331_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1140__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0332_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1130__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0332_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1421__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0333_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1135__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0333_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1801__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1554__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1553__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1134__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1132__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1143__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0335_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1133__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0335_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1144__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0336_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1134__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0336_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1728__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0337_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1135__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0337_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1823__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1820__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1184__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1164__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1145__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1485__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1430__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1428__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1260__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1140__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1475__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1429__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1226__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1213__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1139__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1149__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0341_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1147__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0341_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1140__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0341_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1432__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0342_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1145__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0342_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1801__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1737__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1735__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1582__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1144__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1798__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1736__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1555__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1543__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1143__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1152__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0345_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1150__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0345_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1144__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0345_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1739__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0346_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1145__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0346_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1486__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1477__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1227__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1149__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1147__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1157__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0348_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0348_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1158__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0349_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1149__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0349_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1440__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1153__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1162__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0351_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1151__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0351_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1163__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1152__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1748__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0353_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1153__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0353_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1254__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0354_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1155__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0354_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1476__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1283__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1209__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1199__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1156__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1487__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1445__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1444__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1443__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1158__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1168__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0357_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1166__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0357_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1158__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0357_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1449__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0358_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1164__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0358_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1579__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0359_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1160__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0359_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1791__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1601__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1540__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1533__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1161__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1790__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1752__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1751__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1163__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1172__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0362_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1170__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0362_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1163__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0362_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1757__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0363_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1164__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0363_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1489__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1230__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1208__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1168__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1166__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1177__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0365_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1167__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0365_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1192__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0366_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1178__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0366_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1168__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0366_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1457__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0367_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1173__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0367_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1606__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1559__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1539__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1172__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1170__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1182__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0369_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1171__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0369_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1188__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0370_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1183__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0370_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1172__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0370_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1766__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0371_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1173__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0371_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1249__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0372_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1175__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0372_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1489__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1285__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1234__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1233__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1490__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1461__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1192__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1178__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1192__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0375_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1178__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0375_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1465__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0376_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1184__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0376_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1577__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0377_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1180__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0377_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1796__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1603__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1563__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1562__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1181__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1784__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1771__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1770__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1188__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1183__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1188__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0380_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1183__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0380_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1774__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0381_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1184__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0381_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1563__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0382_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1186__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0382_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1812__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1604__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1565__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1562__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1187__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1813__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1780__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1779__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1778__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1188__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1782__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0385_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1194__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0385_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1234__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0386_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1190__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0386_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1491__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1287__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1236__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1233__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1191__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1492__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1471__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1470__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1469__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1192__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1473__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0389_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1193__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0389_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1194__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0390_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1473__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0391_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1465__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0391_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1449__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0391_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1196__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0391_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1432__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1425__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1414__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1392__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1385__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1332__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1289__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1236__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1234__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1233__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1487__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1435__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1356__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1209__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1199__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1231__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0395_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1252__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0396_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1250__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0396_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1205__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0396_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1487__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1476__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1322__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1205__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1282__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0398_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1257__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0398_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1257__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0398_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1203__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0398_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1487__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1438__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1437__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1434__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1205__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1485__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1365__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1210__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1205__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1231__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0401_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1355__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0402_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1352__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0402_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1207__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0402_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1516__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1475__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1230__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1208__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1230__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0404_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1209__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0404_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1231__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0405_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1511__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1510__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1475__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1361__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1227__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1308__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0407_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1212__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0407_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1508__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1507__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1303__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1226__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1213__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1227__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0409_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1224__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0410_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1215__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0410_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1504__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1503__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1317__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1307__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1225__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1501__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0412_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1500__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0412_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1482__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0412_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1222__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0412_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1498__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1336__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1313__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1221__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1220__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1312__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0414_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1219__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0414_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1498__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1493__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1350__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1337__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1220__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1222__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0416_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1222__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0417_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1225__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0418_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1481__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1394__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1345__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1343__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1224__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1225__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0420_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1226__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0421_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1227__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0422_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1231__A4 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0423_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1297__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0424_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1296__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0424_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1229__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0424_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1486__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1477__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1230__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1231__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0426_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1235__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0427_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1488__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1451__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1325__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1234__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1233__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1235__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0429_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1235__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0430_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1236__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0431_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1412__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0432_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1396__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0432_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1389__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0432_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1237__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0432_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1388__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0433_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1241__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0433_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1240__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0434_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1240__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0435_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1397__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0436_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1241__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0436_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1245__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0437_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1242__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0437_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1243__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0438_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1391__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0439_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1390__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0439_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1244__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0439_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1385__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0440_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1385__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0441_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1375__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0442_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1330__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0442_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1247__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0442_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1526__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1525__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1468__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1376__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1331__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1603__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0444_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1577__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0444_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1285__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0444_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1249__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0444_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1327__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0445_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1285__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0445_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1488__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1456__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1454__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1452__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1284__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1602__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0447_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1578__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0447_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1284__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0447_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1252__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0447_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1290__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0448_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1284__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0448_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1601__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0449_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1579__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0449_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1283__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0449_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1254__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0449_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1292__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0450_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1283__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0450_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1257__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0451_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1256__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0451_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1600__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1580__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1580__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1282__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1257__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1295__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0453_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1295__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0453_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1282__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0453_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1582__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0454_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1260__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0454_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1280__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0455_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1260__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0455_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1299__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0456_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1299__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0456_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1279__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0456_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1417__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0457_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1298__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0457_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1264__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0457_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1264__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0457_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1264__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0458_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1263__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0458_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1633__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1584__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1584__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1298__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1264__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1302__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0460_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1302__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0460_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1298__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0460_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1279__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0460_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1586__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0461_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1267__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0461_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1277__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0462_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1267__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0462_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1306__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0463_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1306__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0463_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1276__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0463_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1304__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0464_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1270__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0464_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1270__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0464_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1615__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1588__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1305__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1270__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1270__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1309__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0466_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1309__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0466_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1305__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0466_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1276__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0466_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1312__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0467_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1274__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0467_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1590__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0468_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1273__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0468_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1313__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0469_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1310__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0469_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1274__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0469_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1314__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0470_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1275__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0470_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1309__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0471_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1309__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0471_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1305__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0471_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1276__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0471_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1278__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0472_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1278__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0473_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1302__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0474_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1302__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0474_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1298__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0474_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1279__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0474_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1281__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0475_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1281__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0476_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1295__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0477_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1295__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0477_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1282__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0477_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1293__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0478_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1293__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0478_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1283__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0478_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1291__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0479_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1284__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0479_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1328__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0480_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1328__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0480_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1285__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0480_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1288__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0481_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1604__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0482_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1287__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0482_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1288__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0483_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1331__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0484_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1330__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0484_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1490__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1489__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1460__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1329__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1326__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1291__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0486_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1325__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0487_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1323__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0487_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1293__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0488_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1293__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0488_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1322__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0489_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1294__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0489_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1321__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0490_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1297__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0491_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1296__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0491_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1321__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0492_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1320__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0493_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1299__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0494_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1299__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0494_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1301__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0495_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1300__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0495_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1320__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0496_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1319__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0497_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1308__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0498_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1303__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0498_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1319__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0499_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1481__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1400__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1398__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1393__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1305__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1306__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0501_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1306__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0501_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1317__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0502_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1307__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0502_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1318__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0503_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1318__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0504_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1316__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0505_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1315__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0505_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1314__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0506_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1312__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0507_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1313__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0508_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1314__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0509_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1316__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0510_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1315__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0510_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1317__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0511_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1317__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0512_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1318__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0513_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1319__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0514_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1320__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0515_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1321__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0516_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1324__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0517_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1323__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0518_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1324__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0519_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1325__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0520_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1329__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0521_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1326__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0521_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1330__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0522_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1328__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0523_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1328__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0523_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1329__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0524_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1330__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0525_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1468__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0526_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1331__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0526_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1407__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0527_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1382__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0527_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1377__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0527_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0528_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1522__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0528_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1333__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0528_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1375__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0529_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1497__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0530_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1480__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0530_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1386__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0530_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1370__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0530_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1338__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0530_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1370__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0531_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1338__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0531_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1338__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0532_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1338__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0533_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1370__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0534_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0534_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1345__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0535_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1343__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0535_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1483__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0536_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1482__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0536_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1408__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0536_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1343__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0536_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1342__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0536_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1672__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0537_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1343__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0537_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1342__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0537_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1371__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0538_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1345__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0538_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1371__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0539_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1344__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0539_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1345__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0540_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1371__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0541_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1367__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0541_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1667__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0542_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1661__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0542_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1363__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0542_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1357__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0542_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1666__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0543_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1365__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0543_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1349__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0543_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1484__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0544_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1478__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0544_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1416__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0544_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1365__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0544_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1349__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0544_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1372__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0545_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1357__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0545_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1357__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0546_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1656__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0547_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1655__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0547_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1356__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0547_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1355__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0547_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1353__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0548_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1373__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0549_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1354__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0549_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1356__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0550_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1373__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0551_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1356__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0551_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1369__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0552_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1357__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0552_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1367__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0553_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1520__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0554_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1519__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0554_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1489__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0554_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1359__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0554_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1360__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0555_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1368__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0556_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1366__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0556_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1373__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0557_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1366__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0557_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1675__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0558_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1667__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0558_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1363__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0558_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1374__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0559_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1366__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0559_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1665__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0560_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1365__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0560_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1372__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0561_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1366__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0561_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1367__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0562_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1375__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0563_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1374__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0564_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1373__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0565_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1371__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0566_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1372__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0567_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1373__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0568_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1374__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0569_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1375__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0570_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1467__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0571_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1376__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0571_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1406__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0572_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1381__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0572_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1377__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0572_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1452__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0573_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1418__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0573_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1378__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0573_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1434__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0574_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1409__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0574_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1393__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0574_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1387__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0574_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1379__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0574_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1385__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0575_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1436__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0576_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1405__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0576_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1395__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0576_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1391__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0576_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1384__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0576_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1451__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0577_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1435__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0577_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1394__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0577_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1386__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0577_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1383__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0577_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1451__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0578_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1435__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0578_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1394__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0578_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1386__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0578_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1383__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0578_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1384__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0579_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1385__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0580_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1392__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0581_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1392__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0582_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1457__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0583_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1440__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0583_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1420__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0583_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1403__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0583_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1389__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0583_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1391__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0584_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1390__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0584_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1392__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0585_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1392__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0586_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1404__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0587_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1395__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0588_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1404__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0589_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1473__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0590_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1465__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0590_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1449__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0590_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1439__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0590_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1401__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0590_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1400__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0591_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1398__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0591_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1411__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0592_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1399__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0592_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1410__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0593_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1400__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0593_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1401__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0594_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1404__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0595_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1474__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0596_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1466__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0596_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1453__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0596_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1440__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0596_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1403__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0596_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1404__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0597_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1527__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0598_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1450__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0598_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1433__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0598_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1426__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0598_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1415__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0598_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1460__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0599_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1442__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0599_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1427__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0599_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1416__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0599_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1408__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0599_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1460__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0600_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1442__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0600_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1427__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0600_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1416__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0600_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1408__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0600_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1415__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0601_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1415__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0602_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1413__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0603_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1424__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0604_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1422__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0604_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1413__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0604_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1472__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0605_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1432__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0605_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1431__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0605_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1414__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0605_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1413__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0605_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1415__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0606_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1415__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0607_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1426__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0608_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1484__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0609_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1478__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0609_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1424__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0609_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1422__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0609_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1419__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0609_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1469__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0610_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1461__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0610_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1443__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0610_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1428__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0610_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1419__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0610_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1426__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0611_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1464__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0612_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1458__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0612_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1448__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0612_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1425__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0612_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1421__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0612_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1426__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0613_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1430__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0614_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1423__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0614_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1429__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0615_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1424__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0615_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1425__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0616_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1426__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0617_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1433__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0618_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1433__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0619_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1431__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0620_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1438__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0621_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1437__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0621_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1431__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0621_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1433__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0622_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1433__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0623_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1441__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0624_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1436__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0625_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1441__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0626_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1445__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0627_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1444__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0627_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1438__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0627_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1439__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0628_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1441__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0629_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1441__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0630_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1450__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0631_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1450__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0632_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1448__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0633_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1446__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0634_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1456__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0635_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1454__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0635_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1447__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0635_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1448__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0636_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1450__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0637_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1450__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0638_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1453__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0639_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1453__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0640_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1459__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0641_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1462__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0642_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1455__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0642_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1463__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0643_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1456__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0643_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1458__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0644_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1458__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0645_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1459__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0646_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1466__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0647_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1466__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0648_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1464__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0649_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1471__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0650_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1470__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0650_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1464__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0650_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1466__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0651_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1466__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0652_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1468__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0653_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1474__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0654_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1474__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0655_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1472__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0656_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1472__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0657_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1474__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0658_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1474__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0659_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1486__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0660_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1487__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0661_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1477__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0661_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1486__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0662_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1485__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0663_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1481__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0664_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1481__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0665_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1483__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0666_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1483__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0667_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1484__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0668_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1485__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0669_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1486__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0670_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1488__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0671_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1488__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0672_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1490__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0673_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1490__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0674_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1491__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0675_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1492__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0676_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1527__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0677_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1526__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0677_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0677_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1493__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0677_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1845__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0678_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1843__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0678_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1505__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0678_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1502__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0678_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1499__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0678_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1524__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0679_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1521__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0679_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1518__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0679_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1515__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0679_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1496__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0679_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1512__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0680_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1509__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0680_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1505__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0680_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1502__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0680_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1499__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0680_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1499__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0681_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1501__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0682_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1500__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0682_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1499__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0682_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1502__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0683_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1504__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0684_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1503__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0684_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1502__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0684_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1508__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0685_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1507__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0685_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1505__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0685_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1505__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0686_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1521__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0687_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1518__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0687_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1515__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0687_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1512__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0687_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1509__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0687_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1509__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0688_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1511__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0689_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1510__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0689_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1509__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0689_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1512__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0690_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1514__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0691_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1513__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0691_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1512__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0691_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1515__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0692_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1517__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0693_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1516__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0693_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1515__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0693_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1520__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0694_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1519__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0694_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1518__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0694_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1518__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0695_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1521__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0696_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1523__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0697_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1522__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0697_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1521__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0697_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1526__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0698_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1525__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0698_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1524__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0698_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1524__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0699_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1526__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0700_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1782__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0701_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1774__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0701_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1757__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0701_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1529__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0701_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1739__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0702_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1732__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0702_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1722__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0702_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1700__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0702_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1693__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0702_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1796__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0703_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0703_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1563__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0703_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1562__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0703_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0703_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1784__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0704_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1769__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0704_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1649__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0704_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1646__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0704_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1565__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0704_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1656__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0705_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1638__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0705_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1557__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0705_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1540__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0705_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1533__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0705_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1560__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0706_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1760__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0707_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1602__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0707_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1578__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0707_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1537__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0707_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1741__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0708_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1600__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0708_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1580__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0708_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1580__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0708_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1537__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0708_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1801__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0709_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0709_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1640__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0709_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1636__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0709_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1537__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0709_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1560__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0710_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1558__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0711_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1539__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0711_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1559__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0712_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1540__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0712_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1560__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0713_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1829__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0714_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1828__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0714_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1798__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0714_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1662__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0714_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1556__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0714_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1801__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0715_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1665__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0715_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1555__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0715_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1543__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0715_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1556__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0716_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1613__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0717_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1554__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0717_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1553__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0717_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1794__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0718_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1788__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0718_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1672__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0718_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1660__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0718_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1551__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0718_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1658__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0719_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1622__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0719_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1550__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0719_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1549__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0719_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1620__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0720_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1619__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0720_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1548__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0720_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1817__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0721_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1814__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0721_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1671__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0721_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1657__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0721_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1549__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0721_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1551__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0722_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1551__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0723_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1554__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0724_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1819__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0725_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1818__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0725_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1702__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0725_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1625__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0725_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1553__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0725_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1554__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0726_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1555__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0727_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1556__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0728_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1560__A4 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0729_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1832__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0730_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1831__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0730_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1559__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0730_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1835__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0731_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1834__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0731_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1655__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0731_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1654__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0731_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1559__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0731_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1560__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0732_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1564__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0733_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1667__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0734_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1644__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0734_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1608__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0734_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1563__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0734_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1562__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0734_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1564__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0735_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1564__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0736_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1565__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0737_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1720__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0738_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1704__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0738_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1697__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0738_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1566__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0738_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0739_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1570__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0739_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1569__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0740_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1569__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0741_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1705__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0742_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1570__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0742_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1574__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0743_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1571__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0743_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1572__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0744_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1699__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0745_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1698__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0745_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1573__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0745_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1693__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0746_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1693__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0747_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1683__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0748_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1650__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0748_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1576__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0748_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1845__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0749_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1813__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0749_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1777__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0749_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1684__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0749_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1651__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0749_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1647__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0750_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1603__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0750_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1606__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0751_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1602__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0751_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1610__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0752_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1601__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0752_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1639__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0753_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1639__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0753_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1600__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0753_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1598__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0754_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1582__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0754_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1634__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0755_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1634__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0755_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1597__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0755_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1632__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0756_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1584__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0756_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1584__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0756_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1633__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0757_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1629__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0757_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1629__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0757_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1597__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0757_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1595__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0758_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1586__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0758_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1616__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0759_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1616__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0759_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1594__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0759_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1708__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0760_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1706__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0760_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1701__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0760_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1615__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0760_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1588__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0760_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1624__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0761_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1589__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0761_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1614__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0762_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1594__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0762_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1622__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0763_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1618__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0763_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1591__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0763_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1623__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0764_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1592__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0764_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1624__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0765_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1593__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0765_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1614__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0766_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1594__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0766_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1596__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0767_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1596__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0768_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1633__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0769_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1629__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0769_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1629__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0769_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1597__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0769_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1599__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0770_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1599__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0771_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1639__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0772_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1639__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0772_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1600__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0772_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1611__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0773_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1611__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0773_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1601__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0773_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1607__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0774_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1602__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0774_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1648__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0775_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1648__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0775_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1603__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0775_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1605__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0776_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1605__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0777_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1651__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0778_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1650__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0778_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1607__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0779_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1645__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0780_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1608__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0780_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1645__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0781_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1791__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0782_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1790__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0782_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1750__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0782_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1642__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0782_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1612__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0782_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1611__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0783_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1611__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0783_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1642__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0784_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1612__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0784_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1645__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0785_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1807__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0786_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1805__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0786_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1678__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0786_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1669__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0786_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1627__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0786_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1624__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0787_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1615__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0787_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1616__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0788_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1616__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0788_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1631__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0789_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1617__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0789_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1627__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0790_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1623__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0791_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1787__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0792_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1621__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0792_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1786__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0793_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1621__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0793_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1622__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0794_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1623__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0795_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1626__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0796_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1625__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0796_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1626__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0797_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1625__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0797_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1627__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0798_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1627__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0799_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1637__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0800_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1821__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0801_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1797__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0801_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1788__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0801_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1716__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0801_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1631__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0801_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1636__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0802_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1630__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0802_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1631__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0803_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1637__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0804_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1802__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0805_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1731__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0805_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1729__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0805_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1726__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0805_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1633__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0805_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1634__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0806_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1634__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0806_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1640__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0807_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1636__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0807_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1825__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0808_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1824__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0808_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1802__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0808_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0808_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1636__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0808_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1637__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0809_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1643__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0810_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1793__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0811_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1791__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0811_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0811_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1642__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0811_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1641__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0811_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1642__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0812_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1641__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0812_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1641__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0813_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1643__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0814_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1643__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0815_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1645__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0816_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1785__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0817_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1784__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0817_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1759__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0817_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1675__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0817_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1645__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0817_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1649__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0818_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1646__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0818_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1650__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0819_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1648__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0820_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1648__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0820_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1649__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0821_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1650__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0822_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1777__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0823_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1651__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0823_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1715__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0824_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0824_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0824_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1843__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0825_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1840__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0825_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1653__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0825_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1683__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0826_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1681__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0827_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1656__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0827_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1680__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0828_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1656__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0828_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1681__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0829_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1674__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0829_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1661__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0830_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1817__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0831_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1795__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0831_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1787__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0831_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1671__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0831_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1659__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0831_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1677__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0832_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1661__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0832_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1678__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0833_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1661__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0833_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1674__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0834_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1663__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0835_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1679__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0836_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1664__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0836_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1666__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0837_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1679__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0838_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1666__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0838_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0839_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1674__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0839_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1682__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0840_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1673__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0840_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1838__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0841_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1837__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0841_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1670__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0841_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1679__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0842_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1670__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0842_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1673__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0843_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1677__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0844_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1673__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0844_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1677__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0845_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1673__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0845_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1674__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0846_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1683__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0847_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1682__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0848_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1679__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0849_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1678__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0850_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1679__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0851_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1681__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0852_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1681__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0853_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1682__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0854_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1683__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0855_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0856_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1684__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0856_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1714__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0857_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1689__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0857_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1685__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0857_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1761__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0858_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1725__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0858_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1686__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0858_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1742__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0859_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1717__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0859_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1701__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0859_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1695__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0859_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1687__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0859_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1693__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0860_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1744__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0861_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1713__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0861_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1703__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0861_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1699__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0861_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1692__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0861_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1759__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0862_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1743__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0862_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1702__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0862_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1694__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0862_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1691__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0862_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1759__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0863_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1743__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0863_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1702__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0863_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1694__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0863_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1691__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0863_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1692__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0864_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1693__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0865_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1700__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0866_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1700__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0867_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1766__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0868_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1748__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0868_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0868_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1711__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0868_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1697__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0868_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1699__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0869_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1698__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0869_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1700__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0870_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1700__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0871_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1712__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0872_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1703__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0873_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1712__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0874_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1782__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0875_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1774__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0875_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1757__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0875_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1747__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0875_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1709__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0875_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1708__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0876_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1706__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0876_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1719__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0877_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1707__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0877_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1718__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0878_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1708__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0878_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1709__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0879_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1712__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0880_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1783__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0881_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1775__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0881_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1762__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0881_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1748__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0881_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1711__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0881_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1712__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0882_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1848__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0883_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1758__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0883_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1740__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0883_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1733__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0883_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1723__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0883_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1769__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0884_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1750__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0884_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1734__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0884_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1724__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0884_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1716__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0884_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1769__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0885_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1750__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0885_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1734__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0885_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1724__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0885_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1716__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0885_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1723__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0886_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1723__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0887_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1721__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0888_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1731__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0889_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1729__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0889_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1721__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0889_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1781__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0890_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1739__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0890_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1738__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0890_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1722__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0890_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1721__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0890_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1723__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0891_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1723__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0892_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1733__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0893_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1778__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0894_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1770__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0894_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1751__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0894_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1735__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0894_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1726__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0894_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1733__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0895_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1773__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0896_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1767__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0896_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1756__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0896_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1732__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0896_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1728__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0896_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1733__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0897_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1737__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0898_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1730__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0898_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1736__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0899_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1731__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0899_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1732__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0900_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1733__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0901_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1740__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0902_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1740__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0903_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1738__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0904_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1746__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0905_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1745__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0905_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1738__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0905_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1740__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0906_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1740__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0907_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1793__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0908_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1791__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0908_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1746__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0908_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1745__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0908_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1742__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0908_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1749__A1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0909_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1744__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0910_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1749__A2_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0911_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1753__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0912_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1752__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0912_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1746__B1_N (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0912_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1747__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0913_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1749__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0914_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1749__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0915_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1758__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0916_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1758__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0917_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1756__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0918_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1754__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0919_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1765__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0920_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1763__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0920_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1755__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0920_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1756__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0921_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1758__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0922_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1921__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0923_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1922__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0924_)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_0_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_0_16_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_0_32_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_0_48_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clk_0_48)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_1_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_0_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_0_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1852__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1853__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1854__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1855__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1856__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1857__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1858__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1859__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1861__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1851__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1860__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1862__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1863__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1864__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1865__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1866__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_0_16_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_0_16_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1867__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1868__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1869__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1870__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1871__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1872__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1873__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1874__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1886__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1887__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1888__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1889__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1890__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1891__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1892__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1893__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_16)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_clk_0_32_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_clk_0_32_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1914__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1915__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1916__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1917__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1918__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1919__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1920__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1894__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1895__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1896__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1897__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1909__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1910__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1911__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1912__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1913__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1__leaf_clk_0_32)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_0_48_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_48)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_0_48_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_0_48)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1923__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_0_48)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1924__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_0_48)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_1_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_1_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__CTS_buf_1_0_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__CTS_buf_1_48_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__CTS_buf_1_16_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_1_0)
);

sky130_fd_sc_hd__diode_2 ANTENNA__CTS_buf_1_32_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_clk_1_0)
);

sky130_fd_sc_hd__decap_4 FILLER_0_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_401 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_463 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_1_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_1_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_1_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_2_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_2_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_2_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_3_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_3_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_5_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_403 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_7_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_7_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_7_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_338 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_7_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_7_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_7_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_7_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_7_464 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_8_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_8_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_8_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_9_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_9_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_9_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_9_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_9_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_401 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_405 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_9_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_9_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_11_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_11_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_11_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_11_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_11_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_399 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_460 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_12_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_12_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_13_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_13_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_13_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_465 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_14_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_14_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_14_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_14_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_403 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_14_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_14_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_15_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_15_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_17_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_17_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_17_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_17_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_17_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_17_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_18_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_18_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_18_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_19_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_338 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_19_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_401 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_405 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_19_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_460 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_431 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_21_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_21_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_21_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_21_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_21_461 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_22_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_22_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_23_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_23_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_23_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_23_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_23_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_23_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_23_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_25_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_25_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_25_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_25_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_25_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_25_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_25_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_431 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_27_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_27_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_27_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_29_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_29_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_29_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_29_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_29_463 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_30_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_30_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_30_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_31_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_31_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_31_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_31_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_31_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_33_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_33_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_33_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_33_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_33_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_33_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_33_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_33_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_33_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_33_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_35_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_35_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_35_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_35_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_35_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_405 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_35_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_465 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_36_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_401 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_38_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_368 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_453 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_39_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_39_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_39_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_39_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_39_460 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_40_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_41_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_41_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_41_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_431 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_43_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_43_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_43_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_44_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_44_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_45_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_45_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_45_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_45_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_45_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_45_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_45_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_45_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_46_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_47_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_47_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_49_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_49_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_50_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_50_403 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_51_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_51_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_51_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_51_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_51_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_52_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_52_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_53_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_53_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_53_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_53_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_53_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_53_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_53_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_54_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_54_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_54_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_54_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_54_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_54_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_54_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_54_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_54_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_54_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_55_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_96 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_55_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_55_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_55_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_55_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_55_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_55_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_55_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_55_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_55_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_55_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_55_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_55_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_56_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_56_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_56_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_56_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_56_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_56_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_56_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_56_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_56_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_56_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_56_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_57_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_57_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_57_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_57_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_57_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_57_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_57_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_57_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_57_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_57_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_57_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_57_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_57_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_57_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_57_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_57_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_57_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_57_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_58_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_58_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_58_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_58_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_58_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_58_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_58_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_58_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_58_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_58_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_58_437 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_58_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_58_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_455 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_58_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_58_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_59_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_59_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_59_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_59_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_59_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_59_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_59_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_59_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_59_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_59_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_59_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_403 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_59_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_59_422 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_59_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_59_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_60_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_60_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_60_390 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_60_414 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_60_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_60_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_60_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_60_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_61_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_61_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_61_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_61_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_61_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_61_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_61_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_61_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_61_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_61_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_61_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_61_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_61_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_61_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_61_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_61_458 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_62_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_62_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_62_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_62_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_62_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_62_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_62_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_62_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_62_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_62_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_62_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_62_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_62_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_62_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_62_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_62_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_62_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_63_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_63_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_63_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_63_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_63_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_63_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_63_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_63_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_63_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_63_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_63_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_63_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_63_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_63_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_63_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_63_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_63_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_63_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_64_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_64_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_64_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_64_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_64_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_64_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_64_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_64_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_64_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_64_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_64_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_64_431 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_64_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_64_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_64_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_64_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_65_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_65_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_65_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_65_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_65_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_65_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_65_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_65_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_65_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_65_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_417 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_65_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_65_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_445 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_65_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_65_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_66_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_66_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_66_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_66_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_66_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_66_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_66_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_368 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_66_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_66_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_66_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_66_413 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_66_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_66_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_66_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_66_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_67_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_67_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_67_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_67_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_67_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_67_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_67_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_67_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_67_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_67_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_67_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_406 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_67_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_423 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_67_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_67_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_67_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_67_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_68_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_68_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_68_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_68_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_68_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_439 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_68_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_68_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_68_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_68_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_68_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_69_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_69_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_69_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_69_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_69_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_69_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_69_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_69_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_69_388 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_69_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_69_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_69_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_69_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_69_436 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_441 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_69_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_69_461 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_69_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_70_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_70_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_70_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_70_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_70_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_70_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_70_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_70_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_70_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_70_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_70_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_405 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_70_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_70_429 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_70_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_70_443 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_452 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_70_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_70_464 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_71_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_71_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_71_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_71_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_71_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_71_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_71_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_71_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_71_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_71_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_71_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_71_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_396 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_420 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_71_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_71_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_440 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_71_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_71_462 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_72_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_72_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_72_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_72_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_72_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_72_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_72_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_72_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_72_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_407 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_72_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_72_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_72_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_73_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_73_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_73_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_73_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_393 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_416 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_73_424 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_73_442 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_73_446 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_73_460 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_73_468 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_74_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_74_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_74_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_74_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_74_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_74_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_74_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_74_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_395 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_74_409 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_74_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_74_427 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_430 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_444 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_448 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_74_456 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_74_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_74_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_75_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_75_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_75_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_75_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_75_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_75_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_75_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_75_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_75_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_75_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_75_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_75_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_75_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_75_392 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_75_400 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_75_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_419 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_75_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_75_454 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_75_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_76_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_76_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_76_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_76_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_76_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_76_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_76_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_76_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_394 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_410 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_76_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_432 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_76_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_76_451 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_76_457 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_76_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_76_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_77_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_77_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_77_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_77_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_77_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_77_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_391 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_411 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_421 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_425 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_77_428 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_434 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_77_438 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_77_449 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_77_461 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_77_469 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_78_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_78_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_78_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_78_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_78_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_78_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_78_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_389 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_78_398 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_78_402 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_78_408 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_418 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_433 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_450 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_78_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_78_467 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_79_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_79_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_79_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_79_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_79_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_79_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_79_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_79_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_397 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_79_404 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_79_412 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_79_415 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_79_426 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_435 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_79_447 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_79_459 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_79_466 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

endmodule
