* NGSPICE file created from CLK_RECOVERY.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 D Q SET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 D Q RESET_B CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B Y VGND VPWR
.ends

.subckt CLK_RECOVERY BB_IN CLK_IN CLK_OUT DATA_OUT RESET_N SCAN_IN[0] SCAN_IN[10]
+ SCAN_IN[11] SCAN_IN[12] SCAN_IN[13] SCAN_IN[14] SCAN_IN[15] SCAN_IN[16] SCAN_IN[17]
+ SCAN_IN[18] SCAN_IN[19] SCAN_IN[1] SCAN_IN[20] SCAN_IN[21] SCAN_IN[2] SCAN_IN[3]
+ SCAN_IN[4] SCAN_IN[5] SCAN_IN[6] SCAN_IN[7] SCAN_IN[8] SCAN_IN[9] VDD VSS
XFILLER_39_277 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_247 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_280 VSS VDD sky130_fd_sc_hd__fill_1
X_CTS_buf_1_16 _CTS_buf_1_32/A _CTS_buf_1_16/X VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_22_188 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1757__A2 _1709_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1518__B _1524_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_317 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_77_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1534__A _1906_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_406 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1693__B2 _1692_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1693__A1 _1529_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_133 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_155 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1709__A _1709_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1748__A2 _1696_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1874__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_321 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1428__B _1419_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_343 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_12 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_328 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1444__A _1443_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_56 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0986__C _0982_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1270_ _1304_/A _1269_/Y _1304_/A _1269_/Y _1270_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_394 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1684__A1 SCAN_IN[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_225 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1619__A _1092_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1739__A2 _1720_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0985_ _0985_/A _0986_/D VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1634__A1_N _1597_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1606_ _1169_/X SCAN_IN[8] _1578_/X _1607_/B VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_59_306 VSS VDD sky130_fd_sc_hd__fill_2
X_1537_ _1760_/A _1609_/A _1741_/A _1734_/A _1537_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1354__A _1354_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1372__B1 _1365_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1468_ _1525_/A _1467_/Y _1468_/C _1468_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1124__B1 _1123_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1399_ _1398_/X _1399_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_27_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1897__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1529__A _1529_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0938__B1 _0937_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_87 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_346 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1363__B1 _1240_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_114 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1666__A1 _1347_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_247 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_269 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1439__A _1401_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1174__A _1463_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_68_125 VSS VDD sky130_fd_sc_hd__fill_2
X_1322_ _1442_/A _1322_/B _1322_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_1_390 VSS VDD sky130_fd_sc_hd__fill_1
X_1253_ SCAN_IN[7] _1579_/B VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1106__B1 _1105_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_342 VSS VDD sky130_fd_sc_hd__fill_2
X_1184_ _1820_/A _1178_/X _1119_/X _1183_/X _1184_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XFILLER_20_423 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1349__A _1347_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0968_ _0968_/A _0968_/B _0968_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1188__A3 _1908_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1068__B _1068_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_28 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1084__A _1084_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1345__B1 _1342_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1515__C _1515_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1812__A _1812_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_180 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1648__B2 _1647_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_375 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_55_353 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_702 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_239 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_735 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_367 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_768 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_445 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1259__A _1259_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1584__B1 _1632_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1912__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1706__B _1706_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_132 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_143 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_9 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_72 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1639__B2 _1599_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_375 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_194 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_64_60 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_64_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_209 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_389 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_22 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1811__A1 _1789_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1169__A _1906_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1871_ _1871_/D _1871_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_50_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1327__B1 _1249_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_412 VSS VDD sky130_fd_sc_hd__decap_4
X_1305_ _1304_/X _1269_/Y _1276_/C _1270_/X _1305_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1632__A _1632_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1236_ _1191_/A _1332_/A _1240_/A _1235_/X _1237_/A VSS VDD sky130_fd_sc_hd__a211o_4
X_1167_ _1166_/X _1167_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_37_353 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_375 VSS VDD sky130_fd_sc_hd__fill_2
X_1098_ _1271_/A _1098_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_12_209 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1802__A1 _1729_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_231 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_60_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_286 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1921__RESET_B RESET_N VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_27 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1030__A2 _1029_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_415 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1542__A _1630_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1899__D _1899_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_353 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_367 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_510 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_85 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_598 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_202 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1717__A _1719_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_452 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1436__B _1436_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1309__B1 _1276_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1452__A _1452_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_117 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_139 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_342 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_364 VSS VDD sky130_fd_sc_hd__fill_2
X_1021_ _1019_/Y _1018_/B _1022_/C VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__1088__A2 _1066_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_345 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_61_175 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_389 VSS VDD sky130_fd_sc_hd__decap_8
X_1923_ BB_IN _1923_/Q RESET_N _1923_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1854_ _1022_/X _0963_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1260__A2 _1258_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1785_ _1763_/A _1759_/A _1786_/B VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0945__B1_N _0931_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_415 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_106 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1362__A SCAN_IN[19] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_448 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1264__A2_N _1263_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_407 VSS VDD sky130_fd_sc_hd__fill_2
X_1219_ _1219_/A _1219_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1079__A2 _1860_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1512__D _1511_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1081__B _1078_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_172 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_186 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1236__C1 _1235_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_337 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1787__B1 _1619_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_32 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1003__A2 _1002_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_98 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1272__A SCAN_IN[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_201 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_466 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1711__B1 _1762_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_85 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_278 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_440 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_51 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_462 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1490__A2 _1460_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_378 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_153 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_95 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_340 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_94 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_23 VSS VDD sky130_fd_sc_hd__decap_8
X_1570_ _1566_/Y _1705_/B _1571_/B VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1447__A _1447_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1166__B _1157_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_293 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1182__A _1772_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1004_ _0953_/X _1004_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1481__A2 _1394_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_337 VSS VDD sky130_fd_sc_hd__fill_2
X_1906_ _1906_/D _1906_/Q _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
X_1837_ _1837_/A _1836_/C _1837_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1768_ _1768_/A _1767_/Y _1906_/D VSS VDD sky130_fd_sc_hd__or2_4
X_1699_ _1698_/A _1697_/X _1703_/A _1699_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_57_201 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1092__A _1092_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_256 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1820__A _1820_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_13_315 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_40_101 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1870__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_145 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1775__A3 _1770_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_392 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_42 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_53 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_223 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1730__A _1730_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_237 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_63_204 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_131 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_31_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_93 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_170 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_156 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_192 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _1546_/Y _1590_/X _1621_/X _1622_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1177__A _1463_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_396 VSS VDD sky130_fd_sc_hd__fill_1
X_1553_ _1120_/Y _1702_/A _1131_/X _1613_/A _1553_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1484_ _1417_/X _1349_/B _1483_/X _1484_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_39_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1640__A _1734_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_19 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_22_145 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1518__C _1520_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1815__A _1694_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_38 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1678__C1 _1677_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1693__A2 _1573_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1550__A _1108_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_20 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_64 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_86 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_178 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1709__B _1709_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_377 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1725__A _1686_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0986__D _0986_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1444__B _1437_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_82 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_373 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1684__A2 _1777_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_215 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1460__A _1460_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_237 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_36_259 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_229 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1619__B _1619_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0984_ _0984_/A _0985_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__0947__A1 _1870_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1__f_clk_0_32_A clkbuf_0_clk_0_32/X VSS VDD sky130_fd_sc_hd__diode_2
X_1605_ _1603_/X _1605_/B _1605_/X VSS VDD sky130_fd_sc_hd__xor2_4
XANTENNA__1616__A2_N _1615_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1635__A _1630_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1536_ _1536_/A _1734_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1357__D1 _1369_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1372__A1 _1349_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1467_ _1375_/X _1467_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_47_19 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1124__A1 _1719_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1398_ _1304_/X _1397_/X _1398_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_27_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_395 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_29 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_454 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_115 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_22 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_119 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0938__A1 _0928_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1545__A _1552_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1363__A1 _1894_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1363__B2 _1346_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_215 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1666__A2 _1630_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_410 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_421 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_270 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_53_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_262 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1439__B _1438_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1051__B1 _1032_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1455__A _1462_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1321_ _1321_/A _1296_/Y _1320_/Y _1321_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_1252_ _1200_/Y _1578_/B _1252_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1106__A1 _1103_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_351 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_384 VSS VDD sky130_fd_sc_hd__fill_2
X_1183_ _1771_/A _1171_/Y _1182_/X _1183_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1190__A _1189_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_398 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_281 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_240 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1290__B1 _1252_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_402 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1349__B _1349_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0967_ _0968_/A _0968_/B _0967_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1042__B1 _1032_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1084__B _1084_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1345__A1 _1394_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_137 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1515__D _1516_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1519_ _1359_/A _1520_/B _1521_/C VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_59_148 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_118 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1812__B _1811_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1864__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_365 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_70_324 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_313 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_218 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_736 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_379 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_70_346 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_769 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_428 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1259__B SCAN_IN[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1584__B2 _1263_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_402 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_177 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_65_129 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_84 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_14 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_140 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_73_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_72 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_61_335 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_387 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_346 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_34 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1811__A2 _1803_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1870_ _1153_/X _1870_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1648__A1_N _1602_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1185__A _1908_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1327__A1 _1463_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1887__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_1304_ _1304_/A _1304_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_69_457 VSS VDD sky130_fd_sc_hd__fill_2
X_1235_ _1231_/X _1233_/X _1234_/X _1235_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_49_181 VSS VDD sky130_fd_sc_hd__fill_2
X_1166_ _1166_/A _1157_/X _1166_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_37_365 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_64_195 VSS VDD sky130_fd_sc_hd__decap_8
X_1097_ _1096_/Y _1097_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1802__A2 _1724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_390 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1095__A _1094_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1823__A _1820_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_438 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_54 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_98 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_143 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_195 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_20 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_500 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_64 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_379 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_511 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_210 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_599 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1006__B1 _1005_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1717__B _1695_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_74 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1309__B2 _1270_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_276 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_78_265 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1452__B _1378_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_71 VSS VDD sky130_fd_sc_hd__fill_2
X_1020_ _0999_/X _1015_/X _1019_/Y _1011_/B _1022_/B VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1088__A3 _1084_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_151 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1493__B1 _1113_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_357 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_195 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_154 VSS VDD sky130_fd_sc_hd__fill_2
X_1922_ _1922_/D _1847_/B RESET_N _1923_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_42_390 VSS VDD sky130_fd_sc_hd__fill_2
X_1853_ _1853_/D _1853_/Q _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1784_ _1763_/A _1759_/A _1771_/A _1769_/A _1789_/A VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_69_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_419 VSS VDD sky130_fd_sc_hd__decap_3
X_1218_ _1218_/A _1219_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1081__C _1081_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_110 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_184 VSS VDD sky130_fd_sc_hd__fill_2
X_1149_ _1147_/A _1139_/X _1148_/Y _1149_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1484__B1 _1483_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1902__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_154 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1236__B1 _1240_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_349 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1787__A1 _1089_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1818__A _1702_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_239 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_44 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_401 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_412 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1711__A1 _1111_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_257 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_30 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1475__B1 _1138_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_357 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1227__B1 _1213_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_330 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_349 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_363 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1728__A _1728_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_62 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_396 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_46 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_272 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1463__A _1463_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1182__B _1170_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1925__CLK CLK_OUT VSS VDD sky130_fd_sc_hd__diode_2
X_1003_ _0963_/Y _1002_/X _0971_/Y _1003_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1466__B1 _1464_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_316 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_154 VSS VDD sky130_fd_sc_hd__decap_6
X_1905_ _1758_/Y _1905_/Q _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1638__A _1638_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1836_ _1833_/A _1834_/Y _1836_/C _1827_/D _1916_/D VSS VDD sky130_fd_sc_hd__and4_4
X_1767_ _1727_/X _1765_/X _1766_/X _1767_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
X_1698_ _1698_/A _1697_/X _1698_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__1903__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_268 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_227 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1820__B _1821_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_419 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1457__B1 _1897_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1209__B1 _1208_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_327 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1548__A _1619_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_371 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_179 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1448__B1 _1421_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_110 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_452 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_72_61 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_71_293 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_282 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_72 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_160 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1621_ SCAN_IN[0] _1619_/X _1620_/X _1621_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1177__B _1166_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1552_ _1552_/A _1702_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1193__A _1833_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1483_ _1116_/X _1342_/A _1481_/X _1482_/X _1483_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_39_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_205 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1640__B _1634_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_441 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_308 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_455 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_10_319 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1611__B1 _1600_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1368__A _1366_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1819_ _1702_/A _1819_/B _1819_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1518__D _1517_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1815__B _1547_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1678__B1 _1660_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1831__A _1557_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1693__A3 _1574_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1550__B _1546_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_411 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_433 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_139 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_117 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1278__A _1276_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1602__B1 _1578_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_190 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_334 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_308 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_67_50 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_352 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_76_341 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1741__A _1741_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1309__A1_N _1276_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1460__B _1408_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_208 VSS VDD sky130_fd_sc_hd__fill_2
X_0983_ _0983_/A _0937_/X _0984_/A VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_12_190 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_3 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0947__A2 _0931_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1357__C1 _1350_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1604_ _1812_/A SCAN_IN[10] _1908_/Q _1286_/Y _1605_/B VSS VDD sky130_fd_sc_hd__o22a_4
X_1535_ _1904_/Q _1741_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1372__A2 _1371_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1466_ _1402_/X _1460_/Y _1461_/X _1464_/X _1465_/X _1466_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1124__A2 _1110_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_352 VSS VDD sky130_fd_sc_hd__fill_2
X_1397_ _1096_/Y _1098_/Y _1397_/C _1397_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_27_249 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_219 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_293 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1915__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_263 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1098__A _1271_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_138 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_10_127 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0938__A2 _0936_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_109 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_67 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1826__A _1813_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_337 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1363__A2 _1675_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_105 VSS VDD sky130_fd_sc_hd__fill_2
X_CTS_buf_1_0 _CTS_buf_1_0/A _CTS_buf_1_0/X VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1561__A _1567_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_363 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_344 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_227 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_355 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_86 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1295__A1_N _1257_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1051__A1 _0991_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1736__A _1736_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_142 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1233__A1_N _1191_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_175 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1320_ _1320_/A _1300_/Y _1319_/Y _1320_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_78_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_116 VSS VDD sky130_fd_sc_hd__decap_6
X_1251_ SCAN_IN[8] _1578_/B VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1471__A _1469_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1182_ _1772_/A _1170_/X _1182_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1106__A2 _1095_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_311 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1801__A1_N _1737_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1814__B1 _1119_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1290__A1 _1165_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_252 VSS VDD sky130_fd_sc_hd__fill_2
X_0966_ _1865_/Q _1866_/Q _0961_/X _0968_/B VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1042__A1 _1040_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1646__A _1769_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1345__A2 _1339_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_105 VSS VDD sky130_fd_sc_hd__decap_8
X_1518_ _1506_/X _1524_/B _1520_/B _1517_/Y _1893_/D VSS VDD sky130_fd_sc_hd__and4_4
X_1449_ _1158_/X _1401_/A _1196_/A _1449_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1381__A _1376_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_726 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_252 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_263 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_11_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_22 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_418 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_167 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_108 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1291__A _1283_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_26 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_311 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_73_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_366 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_84 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_451 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1327__A2 SCAN_IN[9] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_436 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_469 VSS VDD sky130_fd_sc_hd__fill_1
X_1303_ _1212_/X _1302_/Y _1303_/Y VSS VDD sky130_fd_sc_hd__nor2_4
X_1234_ _1189_/Y _1332_/A _1176_/A _1451_/A _1234_/X VSS VDD sky130_fd_sc_hd__o22a_4
X_1165_ _1165_/A _1166_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_174 VSS VDD sky130_fd_sc_hd__fill_1
X_1096_ _1094_/A _1096_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_20_299 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1458__B1_N _1457_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0949_ _0948_/X _1005_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1095__B _1271_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1823__B _1821_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_44 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_174 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_336 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_358 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_501 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_512 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_199 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_578 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_98 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_545 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_277 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1006__A1 _0957_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1006__B2 _0952_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1286__A SCAN_IN[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_86 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_59_62 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_233 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_59_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_8 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_314 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1493__A1 _1219_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_144 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_166 VSS VDD sky130_fd_sc_hd__fill_2
X_1921_ _1921_/D _1847_/A RESET_N _1924_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_42_380 VSS VDD sky130_fd_sc_hd__decap_8
X_1852_ _1852_/D _0964_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1783_ _1762_/A _1777_/X _1778_/X _1781_/Y _1782_/X _1783_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1196__A _1196_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1854__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_428 VSS VDD sky130_fd_sc_hd__decap_3
X_1217_ _1217_/A _1217_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1081__D _1080_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_325 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1484__A1 _1417_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1148_ _1147_/X _1148_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_25_347 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_196 VSS VDD sky130_fd_sc_hd__fill_1
X_1079_ _1874_/Q _1860_/Q _0928_/Y _0991_/A _1081_/C VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1236__A1 _1191_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1787__A2 _1658_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1818__B _1819_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_12 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_56 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1834__A _1558_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_435 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1172__B1 _1171_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_225 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1711__A2 _1696_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_54 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_428 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_141 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_100 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_420 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1475__B2 _1361_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_196 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_31_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_166 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1227__A1 _1147_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1227__B2 _1226_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_320 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_328 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_339 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1877__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XPHY_353 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1728__B _1727_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_397 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_58 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1744__A _1703_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_262 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1463__B _1463_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1163__B1 _1162_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_417 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1852__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_439 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_247 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_152 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_163 VSS VDD sky130_fd_sc_hd__fill_2
X_1002_ _0968_/A _0968_/B _0969_/X _1002_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1466__B2 _1465_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1466__A1 _1402_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1904_ _1749_/X _1904_/Q _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_30_383 VSS VDD sky130_fd_sc_hd__decap_4
X_1835_ _1558_/X _1831_/X _1836_/C VSS VDD sky130_fd_sc_hd__or2_4
X_1766_ _1172_/X _1696_/X _1688_/A _1766_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1697_ _1089_/X _1696_/X _1091_/Y _1566_/A _1697_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1654__A SCAN_IN[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_236 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_239 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_442 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1820__C _1819_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1457__A1 _1168_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_111 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_144 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1209__A1 _1199_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_45 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_89 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_158 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1829__A _1798_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_350 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_232 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1145__B1 _1119_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_247 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_217 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1448__A1 _1444_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_150 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_161 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_383 VSS VDD sky130_fd_sc_hd__decap_12
X_1620_ _1092_/A _1619_/B _1620_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_8_365 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_398 VSS VDD sky130_fd_sc_hd__fill_2
X_1551_ _1718_/A _1794_/B _1549_/X _1550_/X _1551_/X VSS VDD sky130_fd_sc_hd__o22a_4
X_1482_ _1103_/X _1216_/Y _1116_/X _1342_/A _1482_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1193__B _1193_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_453 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_283 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_412 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1611__B2 _1610_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1818_ _1702_/A _1819_/B _1821_/B VSS VDD sky130_fd_sc_hd__and2_4
X_1749_ _1742_/X _1744_/X _1747_/X _1748_/X _1749_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1375__B1 SCAN_IN[21] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1384__A _1384_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1678__A1 SCAN_IN[14] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1831__B _1828_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_206 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_431 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_99 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_43 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1278__B _1278_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1602__A1 _1760_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1602__B2 _1601_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1915__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1294__A _1238_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_37 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1118__B1 _1117_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_386 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1460__C _1408_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1469__A _1469_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0982_ _0980_/A _0979_/X _0980_/Y _1007_/C _0982_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_32_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_66_3 VSS VDD sky130_fd_sc_hd__decap_4
X_1603_ _1181_/A _1577_/B _1577_/X _1602_/X _1603_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1357__B1 _1349_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1534_ _1906_/Q _1760_/A VSS VDD sky130_fd_sc_hd__inv_8
X_1465_ _1178_/X _1401_/A _1196_/A _1465_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_79_180 VSS VDD sky130_fd_sc_hd__fill_2
X_1396_ _1237_/A _1401_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_67_364 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1817__D1 _1820_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_261 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1379__A _1245_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_286 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_46 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1842__A _1842_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_375 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_206 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_98 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_73_389 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_434 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1289__A _1332_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_297 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1051__A2 _1050_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1736__B _1730_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_198 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_83 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1752__A _1753_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1250_ _1200_/Y _1452_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_1_382 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1902__D _1733_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1181_ _1181_/A _1771_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1471__B _1471_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_389 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1814__A1 _1548_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1199__A _1199_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1290__A2 SCAN_IN[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_415 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_459 VSS VDD sky130_fd_sc_hd__decap_8
X_0965_ _1853_/Q _0968_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1042__A2 _1041_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1646__B _1646_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1517_ _1516_/A _1516_/B _1517_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__1662__A SCAN_IN[16] VSS VDD sky130_fd_sc_hd__diode_2
X_1448_ _1444_/X _1447_/Y _1421_/B _1448_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1355__A1_N _1198_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_172 VSS VDD sky130_fd_sc_hd__fill_2
X_1379_ _1245_/A _1379_/B _1379_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_55_367 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_378 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_727 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_359 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_70_337 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_749 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_275 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_23_286 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_408 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1837__A _1837_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1572__A _1571_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1876__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1291__B _1290_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_345 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_164 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_61_326 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_359 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1877__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_242 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1009__C1 _0995_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1747__A _1709_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_441 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_69_426 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1732__B1 _1529_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1302_ _1278_/Y _1264_/X _1278_/Y _1264_/X _1302_/Y VSS VDD sky130_fd_sc_hd__a2bb2oi_4
X_1233_ _1191_/A _1332_/A _1176_/A _1451_/A _1233_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_64_142 VSS VDD sky130_fd_sc_hd__fill_1
X_1164_ _1820_/A _1158_/X _1119_/X _1163_/X _1871_/D VSS VDD sky130_fd_sc_hd__a22oi_4
XFILLER_37_367 VSS VDD sky130_fd_sc_hd__fill_2
X_1095_ _1094_/X _1271_/A _1095_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_37_389 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_337 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_212 VSS VDD sky130_fd_sc_hd__fill_2
X_0948_ _0948_/A _0947_/X _0948_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_20_267 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1657__A SCAN_IN[11] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_clk_0_0_A clkbuf_0_clk_0_0/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1723__B1 _1721_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1823__C _1822_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_312 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_67 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_502 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_223 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_546 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_289 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_238 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1006__A2 _1003_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1567__A _1567_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_32 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_54 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_433 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_201 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_78_223 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_78_256 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_356 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_61_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_367 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1493__A2 _1492_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_337 VSS VDD sky130_fd_sc_hd__fill_2
X_1920_ _1848_/X _1688_/A _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_42_370 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1650__C1 _1649_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1851_ _1851_/D CLK_OUT _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1782_ _1188_/X _1709_/A _1529_/A _1782_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_6_282 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_69_201 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_267 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_245 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_37_120 VSS VDD sky130_fd_sc_hd__fill_2
X_1216_ _1216_/A _1216_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_1_70 VSS VDD sky130_fd_sc_hd__fill_2
X_1147_ _1147_/A _1139_/X _1147_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_25_315 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1484__A2 _1349_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1078_ _1023_/Y _1869_/Q _1015_/X _1867_/Q _1078_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1236__A2 _1332_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1387__A _1097_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_208 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_68 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1834__B _1831_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1172__A1 _1169_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_237 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_29_77 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1629__A2_N _1584_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_432 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_337 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_43 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_310 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_87 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1227__A2 _1361_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_321 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_189 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_354 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1297__A _1228_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_387 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1744__B _1744_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_285 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1163__A1 _1753_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_215 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1760__A _1760_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1892__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1001_ _0982_/X _1001_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_74_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_410 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1910__D _1910_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1466__A2 _1460_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_123 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_145 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1623__C1 _1622_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1903_ _1740_/Y _1903_/Q _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_30_351 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1000__A _0993_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1834_ _1558_/X _1831_/X _1834_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1765_ _1763_/A _1754_/X _1764_/Y _1765_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_1696_ _1566_/Y _1696_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1654__B _1558_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1909__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_281 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1820__D _1820_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1457__A2 _1388_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_167 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1209__A2 _1198_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_57 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1829__B _1824_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_362 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_23 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_78 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1553__A2_N _1702_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_222 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_244 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1145__A1 _1820_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_277 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1145__B2 _1144_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_215 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_451 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_63_229 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1448__A2 _1447_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_41 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_189 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_151 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_140 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_162 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_395 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_195 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1755__A _1754_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1550_ _1108_/X _1546_/Y _1550_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1905__D _1758_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1481_ _1304_/X _1394_/A _1479_/X _1480_/X _1481_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_79_373 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_11_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1078__A1_N _1023_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_410 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_432 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_270 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_251 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_465 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1072__B1 _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1817_ _1658_/X _1548_/X _1107_/X _1819_/B _1820_/D _1910_/D VSS VDD sky130_fd_sc_hd__a2111oi_4
XFILLER_7_80 VSS VDD sky130_fd_sc_hd__fill_2
X_1748_ _1152_/X _1696_/X _1762_/A _1748_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1375__A1 _1333_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1375__B2 _1247_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1384__B _1384_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1679_ _1676_/Y _1669_/X _1678_/X _1663_/X _1665_/X _1679_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
XANTENNA__1867__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1678__A2 _1805_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_284 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_67 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_137 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_159 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1602__A2 _1578_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_347 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_325 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1575__A _1575_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_358 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1294__B _1322_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1118__A1 _1116_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_251 VSS VDD sky130_fd_sc_hd__decap_4
X_0981_ _0981_/A _0975_/X _1007_/C VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1469__B _1419_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1602_ _1760_/A _1578_/B _1578_/X _1601_/X _1602_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_8_174 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_59_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1357__A1 _1240_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1533_ _1161_/A _1638_/A _1533_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1464_ _1462_/X _1471_/B _1421_/B _1464_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_67_332 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_321 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_67_310 VSS VDD sky130_fd_sc_hd__fill_1
X_1395_ _1384_/A _1394_/Y _1395_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_27_207 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_218 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1817__C1 _1819_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_402 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_413 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1293__B1 _1282_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_276 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1379__B _1379_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_298 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_12_36 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1395__A _1384_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1924__RESET_B RESET_N VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_262 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_43 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1284__B1 _1252_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_243 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1036__B1 _1041_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_287 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1899__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_188 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_166 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1752__B _1745_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_129 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_49_310 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_321 VSS VDD sky130_fd_sc_hd__fill_2
X_1180_ _1179_/Y _1181_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_335 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_64_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_64_346 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1275__B1 _1274_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_210 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1814__A2 _1813_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1199__B _1198_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_427 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_276 VSS VDD sky130_fd_sc_hd__fill_2
X_0964_ _0964_/A _0964_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_1_0_0_clk_0_0_A clkbuf_0_clk_0_0/X VSS VDD sky130_fd_sc_hd__diode_2
X_1516_ _1516_/A _1516_/B _1520_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1662__B _1798_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1447_ _1447_/A _1447_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1378_ _1378_/A _1379_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_67_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1905__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XPHY_717 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_232 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_739 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_243 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_11_449 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1837__B _1836_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_147 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_48_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_58_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_173 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_143 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_132 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_20 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_176 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_42 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1257__B1 _1202_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1009__B1 _0991_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0932__A _1870_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1747__B _1747_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1763__A _1763_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1732__A1 _1727_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1301_ _1238_/D _1299_/X _1319_/A VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1913__D _1913_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1232_ _1894_/Q _1451_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_110 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_324 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_49_184 VSS VDD sky130_fd_sc_hd__decap_4
X_1163_ _1753_/A _1151_/Y _1162_/X _1163_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_37_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_357 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_154 VSS VDD sky130_fd_sc_hd__fill_2
X_1094_ _1094_/A _1094_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_60_371 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_224 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_393 VSS VDD sky130_fd_sc_hd__decap_4
X_0947_ _1870_/Q _0931_/X _0932_/X _0947_/X VSS VDD sky130_fd_sc_hd__a21bo_4
XANTENNA__1657__B _1548_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1882__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1673__A _1673_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1723__A1 _1713_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1723__B2 _1722_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1823__D _1820_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_419 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_408 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_324 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1487__B1 _1443_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_379 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_45 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_503 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_228 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1006__A3 _1004_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1567__B _1609_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_11 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1583__A _1583_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_423 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_456 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_78_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_59_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_430 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_335 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_143 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_46_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_113 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_179 VSS VDD sky130_fd_sc_hd__decap_4
X_1850_ _1922_/D _1850_/LO VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__1650__B1 _1646_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1781_ _1720_/X _1781_/B _1780_/Y _1781_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1908__D _1783_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_419 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_441 VSS VDD sky130_fd_sc_hd__fill_2
X_1215_ _1215_/A _1307_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1146_ _1146_/A _1147_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_37_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_165 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_124 VSS VDD sky130_fd_sc_hd__fill_2
X_1077_ _0973_/A _1076_/Y _0940_/A _1061_/A _1081_/A VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_40_308 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1668__A _1567_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1641__B1 _1640_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1387__B _1379_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_25 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_404 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_426 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1172__A2 _1162_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_408 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_89 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_400 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_11 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_349 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_71_444 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_300 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_77 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_99 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_311 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_21 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_344 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1578__A _1760_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1297__B _1297_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_388 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1699__B1 _1703_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1163__A2 _1151_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_121 VSS VDD sky130_fd_sc_hd__fill_1
X_1000_ _0993_/X _1000_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1466__A3 _1461_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_135 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1623__B1 _1591_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1902_ _1733_/Y _1583_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1861__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1293__A1_N _1282_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1833_ _1833_/A _1831_/X _1832_/Y _1827_/D _1833_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1764_ _1763_/X _1764_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1695_ _1091_/Y _1695_/B _1695_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_72_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_411 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_25_135 VSS VDD sky130_fd_sc_hd__decap_6
X_1129_ _1128_/X _1129_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_21_330 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1398__A _1304_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1145__A2 _1140_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_463 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_422 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_444 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_116 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_152 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_64 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_141 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_130 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_352 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_163 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_378 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0940__A _0940_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1480_ _1097_/X _1334_/X _1480_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1771__A _1771_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_385 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_216 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1921__D _1921_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_282 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_403 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_62_296 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1011__A _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1072__B2 _1873_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_171 VSS VDD sky130_fd_sc_hd__fill_1
X_1816_ _1813_/X _1820_/D VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_7_70 VSS VDD sky130_fd_sc_hd__decap_4
X_1747_ _1709_/A _1747_/B _1747_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1375__A2 _1367_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1678_ SCAN_IN[14] _1805_/B _1660_/X _1677_/X _1678_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_26_24 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_455 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_293 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_127 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_193 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1591__A _1092_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_20 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1118__A2 _1105_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0935__A _1873_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_263 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_90 VSS VDD sky130_fd_sc_hd__fill_2
X_0980_ _0980_/A _0979_/X _0980_/Y VSS VDD sky130_fd_sc_hd__nor2_4
X_1601_ _1161_/A _1579_/B _1579_/X _1600_/X _1601_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_8_186 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1357__A2 _1346_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1916__D _1916_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1532_ _1567_/C _1638_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1463_ _1463_/A _1463_/B _1471_/B VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_4_381 VSS VDD sky130_fd_sc_hd__decap_4
X_1394_ _1394_/A _1383_/B _1386_/C _1394_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1817__B1 _1107_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1293__B2 _1292_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_458 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_26 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1676__A _1676_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1395__B _1394_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_307 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_314 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1808__B1 _1800_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_403 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1284__B2 _1283_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1284__A1 _1452_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_55 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1036__A1 _1033_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_156 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_41 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_78_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_68_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_351 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_130 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__CTS_root_A CLK_IN VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_388 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1275__A1 _1094_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_285 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_288 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1857__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1496__A _1524_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0963_ _0963_/A _0962_/X _0963_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_71_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1515_ _1506_/X _1524_/B _1515_/C _1516_/B _1515_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1446_ _1445_/X _1447_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_4_93 VSS VDD sky130_fd_sc_hd__fill_2
X_1377_ _1382_/A _1376_/X _1378_/A VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_55_325 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_303 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_718 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_328 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_729 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_14 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_159 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_44 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_58_185 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_64_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_369 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_188 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_61_339 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1257__B2 _1255_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_98 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_49 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1009__A1 _1000_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0932__B _0931_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1763__B _1754_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1886__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_428 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1732__A2 _1731_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1300_ _1238_/D _1299_/X _1300_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_1_170 VSS VDD sky130_fd_sc_hd__decap_8
X_1231_ _1199_/X _1205_/X _1209_/Y _1227_/Y _1230_/Y _1231_/X VSS VDD sky130_fd_sc_hd__o41a_4
XFILLER_1_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_461 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1584__A1_N _1632_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_174 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_64_122 VSS VDD sky130_fd_sc_hd__decap_12
X_1162_ _1905_/Q _1150_/X _1162_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_49_196 VSS VDD sky130_fd_sc_hd__fill_2
X_1093_ _1091_/Y _1571_/A _1093_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_64_177 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_328 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_350 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_383 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_247 VSS VDD sky130_fd_sc_hd__fill_2
X_0946_ _0946_/A _0948_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_9_292 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1537__A1_N _1760_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1673__B _1670_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1184__B1 _1119_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1723__A2 _1716_/Y VSS VDD sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk_0_32 _CTS_buf_1_32/X clkbuf_0_clk_0_32/X VSS VDD sky130_fd_sc_hd__clkbuf_16
X_1429_ _1138_/X _1423_/Y _1429_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_55_100 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1487__A1 _1434_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1487__B2 _1442_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_58 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_24 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_504 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_236 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1567__C _1567_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_269 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_75_75 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1104__A _1103_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_158 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_136 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0943__A _0943_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_350 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1650__A1 _1575_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_394 VSS VDD sky130_fd_sc_hd__decap_3
X_1780_ _1778_/A _1772_/X _1780_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_24_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_280 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1924__D _1846_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_111 VSS VDD sky130_fd_sc_hd__decap_6
X_1214_ _1214_/A _1215_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_25_306 VSS VDD sky130_fd_sc_hd__fill_2
X_1145_ _1820_/A _1140_/X _1119_/X _1144_/X _1145_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XANTENNA__1014__A _1014_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_188 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_199 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_158 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_147 VSS VDD sky130_fd_sc_hd__fill_2
X_1076_ _1873_/Q _1076_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1641__A1 _1743_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0929_ _1865_/Q _1866_/Q _1867_/Q _0929_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_75_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_280 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_306 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_144 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_23 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_301 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_345 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1578__B _1578_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_44 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_378 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_88 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1918__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1594__A _1594_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1699__A1 _1698_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_409 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_420 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1769__A _1769_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1623__A1 _1694_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1901_ _1901_/D _1585_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_30_331 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_180 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_191 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1919__D _1845_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1832_ _1557_/Y _1828_/X _1832_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1763_ _1763_/A _1754_/X _1763_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1694_ _1694_/A _1694_/B _1694_/C _1694_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_72_209 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_38_453 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_423 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_434 VSS VDD sky130_fd_sc_hd__fill_1
X_1128_ _1127_/X _1117_/X _1128_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1059_ _1032_/X _1057_/Y _1058_/X _1861_/D VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_40_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1398__B _1397_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1918__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_55 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_56_261 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1302__B1 _1278_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1589__A _1589_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_76 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_142 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_131 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_120 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_153 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_164 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_364 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_197 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_357 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0940__B _0940_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1890__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1306__A1_N _1276_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_342 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1771__B _1763_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_206 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_397 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_39_228 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_0 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1499__A _1502_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_448 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1011__B _1011_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_459 VSS VDD sky130_fd_sc_hd__decap_8
X_1815_ _1694_/A _1547_/A _1819_/B VSS VDD sky130_fd_sc_hd__and2_4
X_1746_ _1745_/A _1745_/B _1745_/X _1747_/B VSS VDD sky130_fd_sc_hd__a21boi_4
XANTENNA__1375__A3 _1374_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1677_ _1659_/X _1671_/X _1672_/X _1677_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_26_36 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_53_264 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_404 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1202__A _1146_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_68 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_18 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1591__B SCAN_IN[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_54 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_378 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_261 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0935__B _0934_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_426 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0951__A _0951_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_154 VSS VDD sky130_fd_sc_hd__decap_12
X_1600_ _1741_/A _1256_/X _1580_/X _1599_/Y _1600_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_8_198 VSS VDD sky130_fd_sc_hd__decap_6
X_1531_ _1796_/B _1769_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1462_ _1461_/A _1462_/B _1462_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1393_ _1304_/X _1379_/B _1393_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_67_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_356 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1813__A1_N _1777_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1817__A1 _1658_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1014_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_297 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1865__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1692__A _1703_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1729_ _1729_/A _1719_/X _1730_/A VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_58_312 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_359 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1808__A1 _1804_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1808__B2 _1801_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_23 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1284__A2 _1578_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_426 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_201 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_256 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1036__A2 _1034_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_135 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_179 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_53 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1107__A _1494_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0946__A _0946_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_337 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_370 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1275__A2 SCAN_IN[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_256 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1777__A _1777_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0962_ _0958_/Y _0961_/X _0929_/X _0962_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_32_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1514_ _1513_/A _1511_/X _1516_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_1_1__f_clk_0_16_A clkbuf_0_clk_0_16/X VSS VDD sky130_fd_sc_hd__diode_2
X_1445_ _1443_/A _1437_/X _1445_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1017__A _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_142 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_120 VSS VDD sky130_fd_sc_hd__fill_2
X_1376_ SCAN_IN[21] _1525_/A _1375_/X _1376_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_67_153 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_67_197 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_708 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_201 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_719 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_392 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_245 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1687__A _1571_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_26 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_278 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_138 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_418 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_56 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_73_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_156 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1597__A _1597_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1009__A2 _1008_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_440 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_69_418 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1230_ _1157_/A _1513_/A _1208_/X _1166_/A _1516_/A _1230_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
X_1161_ _1161_/A _1753_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_134 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1855__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1092_ _1092_/A _1571_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_64_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_392 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1300__A _1238_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_215 VSS VDD sky130_fd_sc_hd__fill_2
X_0945_ _1869_/Q _0930_/X _0931_/X _0945_/X VSS VDD sky130_fd_sc_hd__a21bo_4
XFILLER_9_271 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1708__B1 _1707_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1673__C _1671_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1184__B2 _1183_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1184__A1 _1820_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1723__A3 _1717_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1428_ _1430_/A _1419_/B _1428_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_68_451 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_304 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_112 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1487__A2 _1198_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1359_ _1359_/A SCAN_IN[19] _1359_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_28_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_178 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_340 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_505 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_204 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_527 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1210__A _1427_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1567__D _1536_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_77 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_421 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_315 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_348 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_307 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_34_318 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1104__B _1095_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1120__A _1585_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1650__A2 _1605_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_292 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_69_237 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1790__A _1753_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1213_ _1138_/X _1212_/X _1213_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_27_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_292 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_421 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_123 VSS VDD sky130_fd_sc_hd__fill_2
X_1144_ _1737_/A _1133_/Y _1143_/X _1144_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_1_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_95 VSS VDD sky130_fd_sc_hd__fill_2
X_1075_ _1071_/Y _1072_/X _1073_/X _1075_/D _1075_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1014__B _1014_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_362 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_181 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1641__A2 _1639_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_395 VSS VDD sky130_fd_sc_hd__decap_3
X_0928_ _1874_/Q _0928_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_20_49 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_417 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_229 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_68_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_101 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_71_424 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_159 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_302 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_373 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_357 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_56 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_379 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1594__B _1589_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_200 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_60 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_266 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1699__A2 _1697_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_93 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1115__A _1114_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_454 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_402 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_167 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1769__B _1716_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_457 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_340 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_362 VSS VDD sky130_fd_sc_hd__decap_4
X_1900_ _1712_/X _1587_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1623__A2 _1618_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_384 VSS VDD sky130_fd_sc_hd__fill_2
X_1831_ _1557_/Y _1828_/X _1831_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1785__A _1763_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_398 VSS VDD sky130_fd_sc_hd__fill_2
X_1762_ _1762_/A _1762_/B _1762_/C _1768_/A VSS VDD sky130_fd_sc_hd__nor3_4
X_1693_ _1529_/X _1573_/Y _1574_/X _1687_/X _1692_/X _1898_/D VSS VDD sky130_fd_sc_hd__o32ai_4
XFILLER_65_240 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1025__A _1023_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_115 VSS VDD sky130_fd_sc_hd__fill_2
X_1127_ _1127_/A _1127_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_446 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_148 VSS VDD sky130_fd_sc_hd__fill_2
X_1058_ _1058_/A _1037_/Y _1058_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_21_310 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_354 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1695__A _1091_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_203 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_56_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1302__B2 _1264_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_295 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_137 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_72_22 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_143 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_298 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_132 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_121 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_110 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_170 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_154 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_99 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_332 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_165 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_314 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_198 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_398 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_369 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_70 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0949__A _0948_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1526__D1 _1492_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_354 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1475__A1_N _1157_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_1 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1499__B _1502_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_276 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_170 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_192 VSS VDD sky130_fd_sc_hd__fill_1
X_1814_ _1548_/X _1813_/X _1119_/X _1909_/D VSS VDD sky130_fd_sc_hd__o21a_4
X_1745_ _1745_/A _1745_/B _1745_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1676_ _1676_/A _1676_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1746__B1_N _1745_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1908__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_48 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_435 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_184 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_5_339 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1220__B1 _1094_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1591__C _1590_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_67_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_240 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1287__B1 _1885_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_416 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_276 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_298 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_162 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_100 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0951__B _0945_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_133 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_166 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_91 VSS VDD sky130_fd_sc_hd__fill_1
X_1530_ _1569_/B _1796_/B VSS VDD sky130_fd_sc_hd__buf_1
X_1461_ _1461_/A _1419_/B _1461_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1392_ _1196_/X _1386_/X _1387_/Y _1390_/Y _1391_/X _1392_/X VSS VDD sky130_fd_sc_hd__a32o_4
XANTENNA__0970__C1 _0969_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_313 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1817__A2 _1548_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1303__A _1212_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_232 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1022__B _1022_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1450__B1 _1448_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1728_ _1728_/A _1727_/X _1728_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1692__B _1692_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1659_ SCAN_IN[12] _1658_/X _1659_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_58_357 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_379 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_37_36 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1808__A2 _1805_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1880__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_69 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1213__A _1138_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_232 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_438 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_235 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1441__B1 _1439_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_10 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_331 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_78_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_386 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_121 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_154 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_49_379 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_64_327 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1123__A _1718_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1871__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_265 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1777__B _1776_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_0961_ _0959_/Y _0961_/B _0961_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1432__B1 _1196_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_3 VSS VDD sky130_fd_sc_hd__decap_4
X_1513_ _1513_/A _1511_/X _1515_/C VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_4_40 VSS VDD sky130_fd_sc_hd__fill_2
X_1444_ _1443_/A _1437_/X _1444_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1017__B _1014_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1375_ _1333_/X _1367_/X _1374_/Y SCAN_IN[21] _1247_/A _1375_/X VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_67_176 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_165 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1033__A _0946_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_709 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1671__B1 SCAN_IN[11] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1687__B _1695_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1749__A2_N _1744_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1853__D _1853_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_408 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1208__A _1166_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_121 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_68 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_246 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1597__B _1584_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1414__B1 _1196_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0957__A _0957_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_49_132 VSS VDD sky130_fd_sc_hd__fill_2
X_1160_ _1579_/A _1161_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_37_327 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_37_349 VSS VDD sky130_fd_sc_hd__fill_2
X_1091_ _1091_/A _1091_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1895__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_371 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1300__B _1299_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0944_ _0951_/A _1068_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1708__A1 _1587_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1184__A2 _1178_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1028__A _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1673__D _1672_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_430 VSS VDD sky130_fd_sc_hd__decap_3
X_1427_ _1427_/A _1408_/B _1408_/C _1427_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1487__A3 _1476_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1358_ _1894_/Q _1359_/A VSS VDD sky130_fd_sc_hd__inv_8
X_1289_ _1332_/A _1460_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1698__A _1698_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_382 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_506 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_59 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_528 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_396 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_227 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1611__A2_N _1610_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_249 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_58 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_415 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_448 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_89 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_59_452 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_33 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_327 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_338 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_444 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_99 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_105 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_382 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1401__A _1401_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_363 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_24_70 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_253 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_205 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1790__B _1790_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1212_ _1211_/Y _1212_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_77_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_30 VSS VDD sky130_fd_sc_hd__decap_3
X_1143_ _1736_/A _1132_/X _1143_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_52_116 VSS VDD sky130_fd_sc_hd__fill_2
X_1074_ _1015_/X _1867_/Q _1871_/Q _0950_/X _1075_/D VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1014__C _1013_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_330 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1311__A _1271_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0927_ _1085_/A _1494_/A _1065_/A _1494_/A _0927_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1314__C1 _1313_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_293 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_56_455 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_330 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_138 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_69 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_303 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_341 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1221__A _1103_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_171 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_336 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1594__C _1614_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_234 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_289 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_219 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_59_271 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_59_260 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_47_466 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1769__C _1716_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1131__A _1583_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_91 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_355 VSS VDD sky130_fd_sc_hd__fill_2
X_1830_ _1827_/A _1828_/X _1829_/Y _1827_/D _1830_/X VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__1785__B _1759_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1761_ _1763_/A _1686_/A _1762_/C VSS VDD sky130_fd_sc_hd__and2_4
X_1692_ _1703_/A _1692_/B _1692_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_57_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_411 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1025__B _1022_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_252 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_414 VSS VDD sky130_fd_sc_hd__fill_2
X_1126_ _1923_/Q _1827_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_25_127 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1041__A _1041_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1057_ _1041_/A _1057_/B _1057_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_33_193 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1695__B _1695_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_49 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1861__D _1861_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_208 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1216__A _1216_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_13 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_211 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_100 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_45 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_71_277 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_133 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_122 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_111 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_155 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_144 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_166 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_337 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_8_304 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_199 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_311 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1526__C1 _1064_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_366 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1126__A _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0965__A _1853_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_230 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_436 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_2 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_469 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1499__C _1497_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_160 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_428 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1796__A _1181_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_141 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_152 VSS VDD sky130_fd_sc_hd__fill_1
X_1813_ _1777_/A _1812_/Y _1778_/A _1811_/X _1813_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_196 VSS VDD sky130_fd_sc_hd__fill_2
X_1744_ _1703_/A _1744_/B _1744_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_7_62 VSS VDD sky130_fd_sc_hd__fill_2
X_1675_ _1675_/A _1759_/A _1675_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_26_447 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_285 VSS VDD sky130_fd_sc_hd__fill_2
X_1109_ _1108_/X _1090_/X _1110_/A VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_53_233 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_428 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1856__D _1031_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_318 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1220__A1 _1103_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1220__B2 _1219_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_78 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1287__B2 _1286_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_425 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1287__A1 _1191_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_233 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_255 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_82 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_450 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_196 VSS VDD sky130_fd_sc_hd__decap_6
X_1460_ _1460_/A _1408_/B _1408_/C _1460_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__0970__B1 _0963_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1391_ _1243_/X _1390_/B _1384_/A _1391_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_79_196 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_67_336 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_380 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1303__B _1302_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_406 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_417 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_428 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1022__C _1022_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_277 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1450__B2 _1449_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1450__A1 _1405_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1727_ _1696_/X _1727_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1658_ _1546_/Y _1658_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1589_ _1589_/A _1589_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_73_306 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_66_391 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1808__A3 _1807_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1213__B _1212_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_244 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_450 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1441__B2 _1440_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1904__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_343 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0952__B1 _0951_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_303 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1489__A1_N _1166_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_325 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1123__B _1110_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_288 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1777__C _1777_/C VSS VDD sky130_fd_sc_hd__diode_2
X_0960_ _1866_/Q _0961_/B VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1432__A1 _1140_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_91 VSS VDD sky130_fd_sc_hd__fill_2
X_1512_ _1506_/X _1502_/B _1510_/Y _1511_/X _1512_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1443_ _1443_/A _1419_/B _1443_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_4_170 VSS VDD sky130_fd_sc_hd__decap_6
X_1374_ _1368_/Y _1373_/Y _1366_/C _1374_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_55_306 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_67_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_309 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1033__B _1029_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_361 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0954__B1_N _0930_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1671__B2 _1548_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1671__A1 SCAN_IN[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1208__B _1516_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_14 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_133 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_328 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_24 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1111__B1 _1110_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_46 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1597__C _1596_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_269 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1414__A1 _1118_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_453 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_424 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1178__B1 _1177_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_457 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_13_94 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_49_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_188 VSS VDD sky130_fd_sc_hd__fill_1
X_1090_ _1089_/X _1092_/A _1090_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1102__B1 _1095_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0973__A _0973_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_361 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_386 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_375 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_206 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_228 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_251 VSS VDD sky130_fd_sc_hd__fill_2
X_0943_ _0943_/A _0951_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1864__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1708__A2 _1706_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1870__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1028__B _0968_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1426_ _1405_/X _1416_/Y _1419_/X _1421_/Y _1425_/X _1879_/D VSS VDD sky130_fd_sc_hd__o32ai_4
X_1357_ _1240_/B _1346_/Y _1349_/X _1350_/X _1369_/A _1357_/X VSS VDD sky130_fd_sc_hd__a2111o_4
XANTENNA__1044__A _1040_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_147 VSS VDD sky130_fd_sc_hd__decap_3
X_1288_ _1285_/X _1287_/X _1288_/X VSS VDD sky130_fd_sc_hd__xor2_4
XANTENNA__1698__B _1697_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_128 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_394 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_507 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_364 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_518 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1864__D _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1219__A _1219_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_57 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1580__B1 _1741_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_456 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_169 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_320 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1401__B _1400_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1893__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_82 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_276 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1129__A _1128_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0968__A _0968_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1211_ _1239_/A _1211_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_65_412 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1323__B1 _1322_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_445 VSS VDD sky130_fd_sc_hd__decap_12
X_1142_ _1903_/Q _1736_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1799__A _1799_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1073_ _1868_/Q _1019_/Y _1868_/Q _1019_/Y _1073_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_169 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_139 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1311__B SCAN_IN[0] VSS VDD sky130_fd_sc_hd__diode_2
X_0926_ _1923_/Q _1494_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1039__A _1032_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1562__B1 _1181_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_209 VSS VDD sky130_fd_sc_hd__fill_2
X_1409_ _1116_/X _1379_/B _1409_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1314__B1 _1274_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_434 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_125 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_158 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_26 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1502__A _1502_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1859__D _1859_/D VSS VDD sky130_fd_sc_hd__diode_2
XPHY_304 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1221__B _1217_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_326 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_194 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1553__B1 _1131_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_209 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1305__B1 _1276_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_412 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_283 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_434 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_286 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1069__C1 _1068_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1412__A _1237_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_180 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_62_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_70 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_183 VSS VDD sky130_fd_sc_hd__fill_2
X_1760_ _1760_/A _1763_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_30_389 VSS VDD sky130_fd_sc_hd__decap_8
X_1691_ _1547_/A _1694_/B _1694_/C _1692_/B VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_32_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_275 VSS VDD sky130_fd_sc_hd__decap_4
X_1125_ _1113_/X _1118_/X _1119_/X _1124_/X _1125_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XFILLER_38_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_437 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1322__A _1442_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1041__B _1034_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1056_ _1058_/A _1060_/B _1057_/B VSS VDD sky130_fd_sc_hd__xor2_4
XFILLER_18_191 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_367 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1783__B1 _1781_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1889_ _1505_/X _1214_/A _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_0_249 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_56_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_253 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1232__A _1894_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_448 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_234 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_57 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_134 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_123 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_112 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_312 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_101 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_156 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_145 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_167 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1774__B1 _1529_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_50 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_323 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1407__A _1382_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1526__B1 _1525_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1142__A _1903_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_415 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_297 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1499__D _1498_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_267 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0981__A _0981_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_109 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1796__B _1796_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_690 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1812_ _1812_/A _1811_/X _1812_/Y VSS VDD sky130_fd_sc_hd__nor2_4
X_1743_ _1743_/A _1694_/B _1694_/C _1744_/B VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1765__B1 _1764_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1674_ _1674_/A _1661_/X _1676_/A _1673_/Y _1674_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__0927__A1_N _1085_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1108_ _1587_/A _1108_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_53_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_289 VSS VDD sky130_fd_sc_hd__decap_12
X_1039_ _1032_/X _1039_/B _1038_/X _1857_/D VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_13_109 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_16 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_153 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_42_49 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1756__B1 _1727_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1220__A2 _1217_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1872__D _1173_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_46 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_35 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_24 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_220 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1287__A2 SCAN_IN[10] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_415 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_286 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1074__A1_N _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_61 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_407 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_72 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_60 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_9 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_93 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1137__A _1259_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0970__A1 _0964_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1390_ _1243_/X _1390_/B _1390_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_4_396 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_67_304 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0976__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1889__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_348 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_392 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_204 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_226 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_462 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1450__A2 _1442_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1738__B1 _1720_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1726_ _1729_/A _1751_/B _1726_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1047__A _1041_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1657_ SCAN_IN[11] _1548_/X _1657_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1588_ _1587_/Y _1269_/Y _1587_/A SCAN_IN[2] _1589_/A VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_58_304 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_337 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_318 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_407 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1510__A _1361_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1867__D _1125_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1441__A2_N _1436_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_127 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_138 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0952__A1 _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_355 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_134 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1911__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_307 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_359 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_57_392 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_223 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_234 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_71 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_395 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1420__A _1388_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1432__A2 _1412_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_292 VSS VDD sky130_fd_sc_hd__fill_2
X_1511_ _1361_/A _1509_/D _1511_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1442_ _1442_/A _1408_/B _1408_/C _1442_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_67_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_101 VSS VDD sky130_fd_sc_hd__decap_12
X_1373_ _1369_/Y _1361_/X _1372_/Y _1355_/X _1354_/A _1373_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
XFILLER_55_329 VSS VDD sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk_0_0 clkbuf_0_clk_0_0/X _1865_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1656__C1 _1655_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_392 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_237 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1671__A2 _1658_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_281 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_292 VSS VDD sky130_fd_sc_hd__decap_4
X_1709_ _1709_/A _1709_/B _1709_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1505__A _1502_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_145 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1111__A1 _1108_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_237 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1240__A _1240_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1414__A2 _1412_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_403 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_13_62 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1178__A1 _1461_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_421 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_163 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_156 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_318 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1102__A1 _1064_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1102__B2 _1101_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1150__A _1904_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_321 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_384 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_398 VSS VDD sky130_fd_sc_hd__fill_2
X_0942_ _0942_/A _0995_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_13_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_263 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_70_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_296 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1028__C _1019_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1425_ _1421_/B _1424_/X _1196_/X _1425_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_68_443 VSS VDD sky130_fd_sc_hd__fill_2
X_1356_ _1198_/X _1351_/Y _1354_/Y _1355_/X _1369_/A VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_55_115 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1044__B _1034_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1287_ _1191_/A SCAN_IN[10] _1885_/Q _1286_/Y _1287_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_63_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_321 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1060__A _1058_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_508 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_192 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_519 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_376 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_59_14 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_428 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_7 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1580__B2 _1256_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1880__D _1880_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_432 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_79 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_398 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_251 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_450 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0968__B _0968_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_7 VSS VDD sky130_fd_sc_hd__decap_4
X_1210_ _1427_/A _1361_/A VSS VDD sky130_fd_sc_hd__inv_8
X_1141_ _1903_/Q _1737_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1323__A1 _1894_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_457 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0984__A _0984_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_148 VSS VDD sky130_fd_sc_hd__decap_4
X_1072_ _1872_/Q _1040_/X _0976_/A _1873_/Q _1072_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_351 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_362 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1087__B1 _1833_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_354 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_173 VSS VDD sky130_fd_sc_hd__decap_8
X_0925_ _0925_/A _1085_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1039__B _1039_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1562__B2 _1608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1055__A _1054_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1408_ _1342_/A _1408_/B _1408_/C _1408_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1314__A1 _1217_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_446 VSS VDD sky130_fd_sc_hd__decap_3
X_1339_ SCAN_IN[13] _1339_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_71_416 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1078__B1 _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_170 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1502__B _1502_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_305 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_140 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_327 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_48 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_51_184 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_24_398 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1875__D _1875_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1002__B1 _0969_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1553__B2 _1613_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1305__A1 _1304_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1305__B2 _1270_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_402 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_59_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_424 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_94 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_298 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_276 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_62_449 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1860__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_310 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1069__B1 _1067_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_354 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_313 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_51_70 VSS VDD sky130_fd_sc_hd__decap_12
X_1690_ _1690_/A _1694_/C VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_51_92 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_435 VSS VDD sky130_fd_sc_hd__fill_1
X_1124_ _1719_/A _1110_/Y _1123_/X _1124_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_38_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1322__B _1322_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1055_ _1054_/X _1060_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_25_107 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_173 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1783__A1 _1762_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1888_ _1502_/X _1216_/A _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1783__B2 _1782_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1883__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1299__B1 _1279_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1513__A _1513_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_287 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_56_276 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_427 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_438 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_124 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_113 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_151 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_102 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_157 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_146 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_135 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_379 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_328 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_168 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1774__A1 _1183_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0982__C1 _1007_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1526__A1 _1525_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_335 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1423__A _1422_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_405 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_254 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_224 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0981__B _0975_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_4 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_151 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_184 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_195 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_680 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ _1789_/X _1803_/Y _1796_/X _1810_/X _1811_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_30_154 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_691 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1257__A1_N _1202_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_165 VSS VDD sky130_fd_sc_hd__decap_6
X_1742_ _1745_/A _1695_/B _1742_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1765__A1 _1763_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_350 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_53 VSS VDD sky130_fd_sc_hd__fill_2
X_1673_ _1673_/A _1670_/X _1671_/X _1672_/X _1673_/Y VSS VDD sky130_fd_sc_hd__nand4_4
XFILLER_38_210 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1333__A _1333_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_254 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_427 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_276 VSS VDD sky130_fd_sc_hd__fill_2
X_1107_ _1494_/A _1107_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1038_ _0950_/X _1037_/Y _1038_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_41_408 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_28 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_42_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1205__B1 _1434_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1756__A1 _1752_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1508__A _1212_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_349 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1243__A _1243_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_298 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_441 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1418__A _1378_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_364 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0970__A2 _1865_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0976__B _0975_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_187 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1639__A2_N _1599_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_360 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1858__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_213 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0992__A _0992_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1683__B1 SCAN_IN[21] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_257 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_238 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_43_290 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1450__A3 _1443_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1725_ _1686_/A _1751_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1738__A1 _1736_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1656_ _1351_/Y _1638_/A _1654_/Y _1655_/X _1674_/A VSS VDD sky130_fd_sc_hd__a211o_4
X_1587_ _1587_/A _1587_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1047__B _1046_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_349 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_58_316 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1063__A _0927_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_360 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1921__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_27 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1510__B _1509_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1426__B1 _1421_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1883__D _1459_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1238__A _1894_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0952__A2 _0947_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_113 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_378 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_179 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_382 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1665__B1 SCAN_IN[15] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1701__A _1587_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_374 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_72_352 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_401 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_434 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_64_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1148__A _1147_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1510_ _1361_/A _1509_/D _1510_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_4_32 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0987__A _0983_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1441_ _1434_/X _1436_/X _1439_/X _1440_/X _1441_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_65 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_113 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_98 VSS VDD sky130_fd_sc_hd__fill_2
X_1372_ _1349_/X _1371_/X _1365_/X _1372_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1656__B1 _1654_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_382 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_249 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_260 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1058__A _1058_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1708_ _1587_/Y _1706_/B _1707_/Y _1709_/B VSS VDD sky130_fd_sc_hd__a21oi_4
X_1639_ _1580_/X _1599_/Y _1580_/X _1599_/Y _1639_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1073__A1_N _1868_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1505__B _1502_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1647__B1 _1577_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_330 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1111__A2 _1090_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1521__A _1506_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1878__D _1415_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1240__B _1240_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_422 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_41 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1178__A2 _1167_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_142 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_60 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_168 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_64_149 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_93 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1102__A2 _1090_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_300 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1150__B _1143_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_396 VSS VDD sky130_fd_sc_hd__fill_2
X_0941_ _0941_/A _0942_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_20_219 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_231 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_220 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1810__B1 _1789_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_275 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1028__D _1028_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1424_ _1417_/X _1411_/X _1423_/Y _1424_/X VSS VDD sky130_fd_sc_hd__a21o_4
Xclkbuf_0_clk_0_48 _CTS_buf_1_48/X clkbuf_0_clk_0_48/X VSS VDD sky130_fd_sc_hd__clkbuf_16
X_1355_ _1198_/A _1351_/Y _1352_/A SCAN_IN[18] _1355_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_19 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_308 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1629__B1 _1596_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_127 VSS VDD sky130_fd_sc_hd__decap_12
X_1286_ SCAN_IN[10] _1286_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_36_341 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1341__A SCAN_IN[14] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1060__B _1060_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_355 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_509 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_388 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_219 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1801__B1 _1131_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1565__C1 _1564_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_26 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1516__A _1516_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_219 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_422 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1251__A SCAN_IN[8] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1580__A1_N _1741_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_396 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_385 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_193 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_54_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_366 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_267 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_81 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1323__A2 _1291_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1140_ _1430_/A _1129_/Y _1139_/X _1140_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_77_296 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_469 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1161__A _1161_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_99 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_66 VSS VDD sky130_fd_sc_hd__fill_2
X_1071_ _1871_/Q _0950_/X _1070_/X _1071_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_65_80 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_374 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_385 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1087__A1 _1085_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_171 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1039__C _1038_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1336__A _1217_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1407_ _1382_/A _1408_/C VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_68_274 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1314__A2 _1310_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_414 VSS VDD sky130_fd_sc_hd__decap_8
X_1338_ _1334_/X _1335_/Y _1336_/X _1337_/Y _1338_/X VSS VDD sky130_fd_sc_hd__a211o_4
X_1269_ SCAN_IN[2] _1269_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_71_428 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1078__B2 _1867_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1502__C _1500_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_306 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_16 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_152 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_317 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_377 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_38 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_27 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_64 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1891__D _1512_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1246__A _1240_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1002__A1 _0968_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_97 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1305__A2 _1269_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_127 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_62_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_428 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1069__A1 _1872_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_160 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_344 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_130 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_325 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_30_369 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_51_82 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1156__A _1199_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0995__A _0995_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_200 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_90 VSS VDD sky130_fd_sc_hd__fill_2
X_1123_ _1718_/A _1110_/A _1123_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_65_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_428 VSS VDD sky130_fd_sc_hd__decap_6
X_1054_ _0991_/A _1045_/X _1054_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_25_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_152 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_336 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_358 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1783__A2 _1777_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1887_ _1499_/X _1217_/A _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_0_218 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1066__A _1084_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_200 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_425 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1299__B2 _1298_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_49 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1513__B _1511_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_469 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_71_269 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_125 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_114 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_450 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_103 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_158 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_147 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_136 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1886__D _1886_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_369 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_169 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1883__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1774__A2 _1709_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0982__B1 _0980_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1526__A2 _1524_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1704__A _1566_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_211 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_93 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_5 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1224__A2_N _1394_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_409 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_174 VSS VDD sky130_fd_sc_hd__fill_2
X_1810_ _1786_/B _1809_/X _1789_/A _1810_/X VSS VDD sky130_fd_sc_hd__o21a_4
XPHY_670 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_122 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_133 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_144 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_692 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1741_ _1741_/A _1745_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1765__A2 _1754_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_373 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_76 VSS VDD sky130_fd_sc_hd__fill_2
X_1672_ _1341_/Y _1544_/A SCAN_IN[13] _1794_/B _1672_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1614__A _1614_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1333__B SCAN_IN[20] VSS VDD sky130_fd_sc_hd__diode_2
X_1106_ _1103_/X _1095_/X _1105_/Y _1106_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_53_225 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_269 VSS VDD sky130_fd_sc_hd__fill_2
X_1037_ _1013_/B _1082_/D _1037_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_21_166 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1205__B2 _1427_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1756__A2 _1755_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1508__B _1503_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1524__A _1100_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1302__A1_N _1278_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_328 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_67_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_255 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_203 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_247 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_280 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_111 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_144 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_137 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_32_73 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_306 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_317 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1434__A _1434_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0992__B _0990_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_225 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1683__B2 _1575_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1683__A1 _1653_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1898__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_91 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_280 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1738__A2 _1745_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1724_ _1724_/A _1716_/B _1716_/C _1724_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1609__A _1609_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1873__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_181 VSS VDD sky130_fd_sc_hd__fill_2
X_1655_ _1351_/Y _1567_/C SCAN_IN[18] _1558_/X _1655_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1586_ _1120_/Y _1265_/Y _1585_/X _1594_/A VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_58_328 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1371__B1 _1343_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1344__A _1343_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1063__B _1063_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_258 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1426__A1 _1405_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_239 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_442 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1426__B2 _1425_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_118 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1519__A _1359_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1238__B _1238_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_14 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_49_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1254__A _1155_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_339 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_169 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_203 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_62 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1665__B2 _1543_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1701__B _1695_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_84 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1920__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1896__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_413 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_453 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1429__A _1138_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1440_ _1149_/X _1388_/X _1402_/X _1440_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_4_44 VSS VDD sky130_fd_sc_hd__fill_2
X_1371_ _1370_/X _1345_/X _1343_/X _1342_/X _1371_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_4_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_67_169 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1656__A1 _1351_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_364 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1339__A SCAN_IN[13] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1058__B _1037_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1707_ _1706_/X _1707_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1592__B1 _1591_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1638_ _1638_/A _1743_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_48_28 VSS VDD sky130_fd_sc_hd__decap_3
X_1569_ _1575_/A _1569_/B _1569_/C _1568_/X _1705_/B VSS VDD sky130_fd_sc_hd__nor4_4
XFILLER_58_125 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1505__C _1503_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_350 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_16 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1647__A1 _1772_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_394 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1521__B _1524_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1240__C _1240_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1894__D _1521_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1249__A _1175_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_434 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_136 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_320 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1102__A3 _1093_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_367 VSS VDD sky130_fd_sc_hd__fill_2
X_0940_ _0940_/A _0940_/B _0941_/A VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1810__A1 _1786_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1159__A _1905_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0998__A _0998_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1911__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk_0_16 _CTS_buf_1_16/X clkbuf_0_clk_0_16/X VSS VDD sky130_fd_sc_hd__clkbuf_16
X_1423_ _1422_/X _1423_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_48_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1354_ _1354_/A _1354_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_68_467 VSS VDD sky130_fd_sc_hd__decap_3
X_1285_ _1176_/A _1577_/B _1249_/X _1284_/X _1285_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_55_139 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1629__B2 _1584_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_353 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_386 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1060__C _1037_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_367 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1801__B2 _1543_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1565__B1 _1575_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_419 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1516__B _1516_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_412 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1317__B1 _1315_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_456 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_37 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_448 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1532__A _1567_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1889__D _1505_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_364 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1562__A2_N _1796_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_24_41 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_24_74 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_257 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1707__A _1706_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1556__B1 _1543_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_73 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_77_231 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_71 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_404 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1442__A _1442_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_320 VSS VDD sky130_fd_sc_hd__decap_12
X_1070_ _1870_/Q _1068_/B _1070_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1087__A2 CLK_OUT VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_150 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_334 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1072__A1_N _1872_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_186 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1617__A _1616_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1336__B SCAN_IN[12] VSS VDD sky130_fd_sc_hd__diode_2
X_1406_ _1376_/X _1408_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_29_19 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_404 VSS VDD sky130_fd_sc_hd__decap_3
X_1337_ SCAN_IN[11] _1219_/X _1337_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1352__A _1352_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1268_ _1268_/A _1304_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_56_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1655__A1_N _1351_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1199_ _1199_/A _1198_/X _1199_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_24_301 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1502__D _1501_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_307 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_323 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_24_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_120 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_318 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_175 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_227 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_238 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1002__A2 _0968_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_201 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_19_117 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1262__A SCAN_IN[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1069__A2 _1040_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_172 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_378 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_95 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_50 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1437__A _1434_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_271 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0995__B _0995_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1122_ _1585_/A _1718_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_256 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_407 VSS VDD sky130_fd_sc_hd__decap_4
X_1053_ _0940_/A _1058_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_18_183 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_194 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_315 VSS VDD sky130_fd_sc_hd__fill_2
X_1886_ _1886_/D _1218_/A _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1783__A3 _1778_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1347__A SCAN_IN[15] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1066__B CLK_OUT VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_17 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1082__A _1082_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_404 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_418 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_115 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_104 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_131 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_148 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_137 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_126 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_159 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_308 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_197 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_370 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0982__A1 _0980_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_42 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_304 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_223 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_47_234 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_278 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1720__A _1566_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_237 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_6 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_120 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_671 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_660 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VSS VDD sky130_fd_sc_hd__fill_2
X_1740_ _1713_/X _1734_/Y _1735_/X _1738_/Y _1739_/X _1740_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1167__A _1166_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_66 VSS VDD sky130_fd_sc_hd__fill_2
X_1671_ SCAN_IN[12] _1658_/X SCAN_IN[11] _1548_/X _1671_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_7_99 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1614__B _1589_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_289 VSS VDD sky130_fd_sc_hd__fill_2
X_1105_ _1104_/X _1105_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1630__A _1630_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1036_ _1033_/X _1034_/X _1041_/A _1039_/B VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_34_451 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_292 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_123 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_178 VSS VDD sky130_fd_sc_hd__decap_4
X_1869_ _1145_/Y _1869_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1805__A _1718_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1524__B _1524_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_245 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1897__D _1527_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_101 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_64 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_410 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_454 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_149 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_85 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1715__A _1690_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_388 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_156 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1434__B _1379_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_82 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1683__A2 _1674_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_440 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_81 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_421 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_3 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_490 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1713_/X _1716_/Y _1717_/X _1721_/Y _1722_/X _1901_/D VSS VDD sky130_fd_sc_hd__o32ai_4
X_1654_ SCAN_IN[18] _1558_/X _1654_/Y VSS VDD sky130_fd_sc_hd__nor2_4
X_1585_ _1585_/A SCAN_IN[3] _1585_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1371__B2 _1342_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1371__A1 _1370_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1063__C _1062_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1270__A2_N _1269_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_215 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1360__A _1359_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_410 VSS VDD sky130_fd_sc_hd__decap_12
X_1019_ _0963_/A _1019_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1426__A2 _1416_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1519__B _1520_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1238__C _1198_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_26 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1535__A _1904_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_303 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1254__B _1579_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_259 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_465 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_51 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1429__B _1423_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_CTS_root CLK_IN _CTS_root/X VSS VDD sky130_fd_sc_hd__clkbuf_16
XANTENNA__1445__A _1443_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_185 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_23 VSS VDD sky130_fd_sc_hd__fill_2
X_1370_ _1334_/X _1335_/Y _1338_/X _1370_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_75_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1180__A _1179_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1656__A2 _1638_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_343 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_284 VSS VDD sky130_fd_sc_hd__fill_2
X_1706_ _1587_/Y _1706_/B _1706_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1592__A1 _1091_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1637_ _1627_/X _1631_/Y _1636_/Y _1637_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1649__B1_N _1648_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1568_ _1630_/A _1544_/A _1552_/A _1694_/A _1568_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_48_18 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1505__D _1504_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1499_ _1502_/A _1502_/B _1497_/X _1498_/X _1499_/X VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__1090__A _1089_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1647__A2 SCAN_IN[9] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1521__C _1521_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_398 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1240__D _1239_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1280__B1 _1259_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1249__B _1577_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1265__A SCAN_IN[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_111 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_148 VSS VDD sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_clk_0_32 clkbuf_0_clk_0_32/X _1911_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_16
XANTENNA__1863__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_310 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_140 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_57_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_162 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_365 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_346 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_200 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1810__A2 _1809_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_255 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_82 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_299 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1175__A _1175_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1422_ _1417_/X _1411_/X _1422_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_68_435 VSS VDD sky130_fd_sc_hd__fill_2
X_1353_ _1352_/X _1354_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_68_457 VSS VDD sky130_fd_sc_hd__fill_1
X_1284_ _1452_/A _1578_/B _1252_/X _1283_/X _1284_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_63_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_365 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_63_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_346 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_398 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_19 VSS VDD sky130_fd_sc_hd__decap_12
X_0999_ _0964_/Y _0999_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1565__A1 _1812_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1085__A _1085_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1317__B2 _1316_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1317__A1 _1307_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1886__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_427 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_118 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_140 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_376 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_346 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_53 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_10_243 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_86 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_203 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1866__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_298 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1556__A1 _1904_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1556__B2 _1555_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_50 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1442__B _1408_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_35 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_37_107 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_460 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_398 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1492__B1 _1491_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_5_280 VSS VDD sky130_fd_sc_hd__decap_3
X_1405_ _1384_/A _1405_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_68_265 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_68_243 VSS VDD sky130_fd_sc_hd__fill_2
X_1336_ _1217_/Y SCAN_IN[12] _1336_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_68_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1352__B SCAN_IN[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_129 VSS VDD sky130_fd_sc_hd__decap_12
X_1267_ _1115_/Y _1265_/Y _1266_/X _1276_/A VSS VDD sky130_fd_sc_hd__o21ai_4
X_1198_ _1198_/A _1198_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_36_140 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_313 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1483__B1 _1481_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_308 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_132 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1235__B1 _1234_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0994__C1 _0993_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_11 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_221 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1543__A _1736_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_53 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_416 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_438 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_246 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_224 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1474__B1 _1472_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_52 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1901__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_452 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_74 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_176 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_187 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1226__B1 _1225_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1718__A _1718_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1437__B _1430_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1453__A _1402_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0995__C _0986_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_70 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_427 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_438 VSS VDD sky130_fd_sc_hd__fill_2
X_1121_ _1120_/Y _1719_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_38_449 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_419 VSS VDD sky130_fd_sc_hd__fill_2
X_1052_ _0991_/A _1050_/X _1051_/Y _1860_/D VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_18_140 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1465__B1 _1196_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_290 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_198 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1628__A _1544_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1885_ _1474_/Y _1885_/Q _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_56_29 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1082__B _1075_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1319_ _1319_/A _1303_/Y _1318_/Y _1319_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1924__CLK _1924_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_238 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1456__B1 _1463_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_116 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_105 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_430 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_24_143 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_149 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_138 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_127 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_316 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_24_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1538__A _1609_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0982__A2 _0979_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1914__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_84 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_7 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_143 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_661 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_371 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_364 VSS VDD sky130_fd_sc_hd__fill_2
X_1670_ SCAN_IN[19] _1837_/A _1669_/X _1670_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_7_397 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_23_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_460 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_408 VSS VDD sky130_fd_sc_hd__fill_2
X_1104_ _1103_/X _1095_/X _1104_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1630__B _1629_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_238 VSS VDD sky130_fd_sc_hd__fill_2
X_1035_ _1011_/B _1041_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_61_260 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1358__A _1894_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1610__B1 _1579_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1868_ _1135_/X _1868_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
X_1799_ _1799_/A _1800_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1805__B _1805_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1093__A _1091_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_39 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1524__C _1524_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_224 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1677__B1 _1672_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1821__A _1716_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_419 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_43 VSS VDD sky130_fd_sc_hd__decap_12
Xclkbuf_0_clk_0_0 _CTS_buf_1_0/X clkbuf_0_clk_0_0/X VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_8_117 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1268__A _1268_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_64 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1601__B1 _1579_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_168 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_57_72 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1683__A3 _1682_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_249 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_208 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_444 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_480 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1124_/X _1720_/X _1529_/X _1722_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_11_190 VSS VDD sky130_fd_sc_hd__fill_1
X_1653_ SCAN_IN[20] _1652_/Y _1653_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1584_ _1632_/A _1263_/X _1632_/A _1263_/X _1584_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1356__C1 _1355_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_308 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1371__A2 _1345_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1018_ _1014_/A _1018_/B _1017_/Y _1853_/D VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_22_422 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1426__A3 _1419_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1238__D _1238_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1816__A _1813_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_359 VSS VDD sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk_0_32 clkbuf_0_clk_0_32/X _1920_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_57_330 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_20 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_396 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_75 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_366 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_274 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1726__A _1729_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1338__C1 _1337_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1445__B _1437_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_197 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_68_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_138 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_116 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1461__A _1461_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_330 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_396 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_75_193 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1813__B1 _1778_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_296 VSS VDD sky130_fd_sc_hd__fill_1
X_1705_ _1093_/X _1705_/B _1706_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1592__A2 SCAN_IN[1] VSS VDD sky130_fd_sc_hd__diode_2
X_1636_ _1734_/A _1634_/X _1724_/A _1629_/X _1636_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
X_1567_ _1567_/A _1609_/A _1567_/C _1536_/A _1569_/C VSS VDD sky130_fd_sc_hd__or4_4
X_1498_ _1217_/Y _1219_/X _1498_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_54_311 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1090__B _1092_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_322 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1521__D _1523_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1280__B2 SCAN_IN[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1280__A1 _1127_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1546__A _1694_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_123 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_1_167 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_77_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_178 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_77_469 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1281__A _1279_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_344 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_62_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_440 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_462 VSS VDD sky130_fd_sc_hd__decap_8
X_1421_ _1130_/X _1421_/B _1421_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_68_447 VSS VDD sky130_fd_sc_hd__fill_2
X_1352_ _1352_/A SCAN_IN[18] _1352_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1283_ _1199_/A _1579_/B _1254_/X _1282_/X _1283_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1191__A _1191_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_322 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_182 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1299__A2_N _1298_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_377 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_314 VSS VDD sky130_fd_sc_hd__fill_1
X_0998_ _0998_/A _1014_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1366__A _1366_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1851__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1565__A2 _1769_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1619_ _1092_/A _1619_/B _1619_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1085__B _1084_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_403 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1317__A2 _1306_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_28 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_333 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_171 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1486__D1 _1485_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_303 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_65 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_215 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1276__A _1276_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1556__A2 _1798_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_95 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_77_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_417 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1442__C _1408_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_72 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_122 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1492__A1 _1469_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_314 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_144 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_358 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_391 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1186__A _1186_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_211 VSS VDD sky130_fd_sc_hd__decap_3
X_1404_ _1393_/X _1395_/X _1401_/X _1403_/X _1404_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1335_ SCAN_IN[12] _1335_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1266_ _1114_/A SCAN_IN[3] _1266_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1197_ _1240_/B _1332_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_36_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1872__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_196 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1483__B2 _1482_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1483__A1 _1116_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_144 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_309 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1235__A1 _1231_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0994__B1 _0991_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1096__A _1094_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_207 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1853__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_56 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1824__A _1724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_233 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1543__B _1543_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_21 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_258 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_314 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1474__B2 _1473_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1474__A1 _1402_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_358 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_464 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1226__A1 _1138_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1718__B _1707_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1734__A _1734_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_251 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1453__B _1451_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0995__D _0995_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1120_ _1585_/A _1120_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_38_406 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_93 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_82 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_65_236 VSS VDD sky130_fd_sc_hd__fill_2
X_1051_ _0991_/A _1050_/X _1032_/X _1051_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_18_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_450 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_61_420 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1465__A1 _1178_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_442 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1876__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1884_ _1466_/Y _1463_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1644__A _1608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1082__C _1081_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1153__B1 _1107_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_428 VSS VDD sky130_fd_sc_hd__decap_3
X_1318_ _1307_/X _1308_/X _1317_/X _1318_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_1249_ _1175_/A _1577_/B _1249_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_64_280 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1456__A1 _1452_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_442 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_106 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_139 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_128 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_117 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_328 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1819__A _1702_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_394 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_66 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1392__B1 _1390_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1144__B1 _1143_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_228 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1899__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XPHY_8 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_261 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_70_294 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_662 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_125 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_695 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1729__A _1729_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_684 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_354 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_372 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_361 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1135__B1 _1107_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_3 VSS VDD sky130_fd_sc_hd__decap_3
X_1103_ _1268_/A _1103_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_53_217 VSS VDD sky130_fd_sc_hd__fill_2
X_1034_ _0950_/X _1028_/X _1034_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1438__A1 _1434_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1843__D1 _1820_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_158 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1610__A1 _1905_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1867_ _1125_/Y _1867_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
X_1798_ _1736_/A _1798_/B _1799_/A VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1374__B1 _1366_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1093__B _1571_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1524__D _1524_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_236 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1677__A1 _1659_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1821__B _1821_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_261 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_55 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_158 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_32 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1601__A1 _1161_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1601__B2 _1600_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_191 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1365__B1 _1347_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_125 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_57_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_51 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_280 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_412 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_294 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1459__A _1453_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_470 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1718_/X _1719_/X _1720_/X _1721_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_7_184 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_7_173 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_162 VSS VDD sky130_fd_sc_hd__decap_4
X_1652_ _1796_/B _1652_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1914__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_1583_ _1583_/A _1632_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1356__B1 _1354_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_228 VSS VDD sky130_fd_sc_hd__fill_2
X_1017_ _1015_/X _1014_/B _1017_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_22_445 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1369__A _1369_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1919_ _1845_/Y _1575_/A _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1595__B1 _1585_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1832__A _1557_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_386 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_389 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_261 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_294 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_405 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1279__A _1279_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1586__B1 _1585_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1726__B _1751_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_132 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1338__B1 _1336_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1742__A _1745_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_371 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1461__B _1419_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_393 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_353 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_161 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_367 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1813__B2 _1811_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1189__A _1885_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1704_ _1566_/A _1709_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1635_ _1630_/A _1724_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1566_ _1566_/A _1566_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1497_ _1334_/X _1218_/A _1497_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1652__A _1796_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_109 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_389 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1099__A _1098_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_426 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1280__A2 SCAN_IN[4] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_448 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_45 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1827__A _1827_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_135 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0__f_clk_0_32_A clkbuf_0_clk_0_32/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_415 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1740__B1 _1738_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_117 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1281__B _1281_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_120 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_52 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_253 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_235 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1008__C1 _1007_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1737__A _1737_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1559__B1 _1169_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1420_ _1388_/X _1421_/B VSS VDD sky130_fd_sc_hd__buf_1
X_1351_ SCAN_IN[17] _1351_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1731__B1 _1730_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1472__A _1412_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_459 VSS VDD sky130_fd_sc_hd__decap_8
X_1282_ _1202_/Y _1256_/X _1257_/X _1281_/Y _1282_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_63_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_345 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_326 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_359 VSS VDD sky130_fd_sc_hd__decap_3
X_0997_ _0996_/X _0998_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1366__B _1361_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1618_ _1590_/X _1618_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1891__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1549_ _1587_/A _1546_/Y _1089_/X _1548_/X _1549_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1722__B1 _1529_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1382__A _1382_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1486__C1 _1477_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_359 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_370 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_392 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_267 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1557__A _1638_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_227 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_32 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1276__B _1270_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_65 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_77_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_84 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_62 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_131 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1492__A2 _1240_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_326 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_348 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_381 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1467__A _1375_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1905__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_271 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_260 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_293 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_201 VSS VDD sky130_fd_sc_hd__decap_8
X_1403_ _1106_/X _1388_/X _1402_/X _1403_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_68_223 VSS VDD sky130_fd_sc_hd__decap_12
X_1334_ _1217_/A _1334_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1265_ SCAN_IN[3] _1265_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_36_120 VSS VDD sky130_fd_sc_hd__decap_4
X_1196_ _1196_/A _1196_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_24_326 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1483__A2 _1342_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_167 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1235__A2 _1233_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_381 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0994__A1 _1061_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1377__A _1382_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1824__B _1822_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1840__A _1652_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_440 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1474__A2 _1468_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_443 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_348 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1226__A2 _1212_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0979__B1_N _0933_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1734__B _1716_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1453__C _1453_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_296 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_76_61 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_204 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1750__A _1790_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_7 VSS VDD sky130_fd_sc_hd__decap_3
X_1050_ _1041_/A _1045_/X _1050_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1900__D _1712_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_270 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1465__A2 _1401_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_134 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_167 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_370 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_392 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_189 VSS VDD sky130_fd_sc_hd__fill_2
X_1883_ _1459_/X _1165_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1197__A _1240_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_204 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1153__B2 _1152_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1153__A1 _1827_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_215 VSS VDD sky130_fd_sc_hd__decap_12
X_1317_ _1307_/A _1306_/Y _1315_/Y _1316_/Y _1317_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_2_80 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1082__D _1082_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1660__A SCAN_IN[13] VSS VDD sky130_fd_sc_hd__diode_2
X_1248_ SCAN_IN[9] _1577_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_71_229 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_207 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1456__A2 _1447_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_462 VSS VDD sky130_fd_sc_hd__decap_8
X_1179_ _1772_/A _1179_/Y VSS VDD sky130_fd_sc_hd__inv_8
XPHY_107 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_129 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_118 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_454 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1819__B _1819_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_362 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1835__A _1558_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1392__A1 _1196_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1392__B2 _1391_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1144__A1 _1737_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1570__A _1566_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_410 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_64 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_292 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_9 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_70_273 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_652 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_137 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_696 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1729__B _1719_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_674 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1923__RESET_B RESET_N VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_351 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1080__B1 _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1745__A _1745_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_377 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1135__B2 _1728_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1135__A1 _1827_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_215 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_237 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1480__A _1097_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1102_ _1064_/X _1090_/X _1093_/X _1095_/X _1101_/X _1102_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
XFILLER_19_440 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_259 VSS VDD sky130_fd_sc_hd__decap_12
X_1033_ _0946_/A _1029_/Y _1033_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1438__A2 _1430_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_421 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_251 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1843__C1 _1844_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_284 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1071__B1 _1070_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1610__A2 SCAN_IN[7] VSS VDD sky130_fd_sc_hd__diode_2
X_1866_ _1112_/X _1866_/Q _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
X_1797_ _1719_/A _1716_/A _1794_/X _1795_/X _1796_/X _1797_/X VSS VDD sky130_fd_sc_hd__a2111o_4
XANTENNA__1374__A1 _1368_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_340 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1390__A _1243_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1677__A2 _1671_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_207 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_410 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_454 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_22 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_44 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1601__A2 _1579_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_77 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_4_369 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1365__A1 _1427_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1365__B2 _1349_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_137 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_321 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_310 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1866__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_229 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_410 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_292 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_95 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_262 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1459__B _1458_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_460 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _1566_/A _1720_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1651_ _1777_/A _1605_/X _1777_/C _1690_/A VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_7_196 VSS VDD sky130_fd_sc_hd__decap_4
X_1582_ _1737_/A _1258_/Y _1581_/X _1597_/A VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1356__A1 _1198_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_398 VSS VDD sky130_fd_sc_hd__fill_2
X_1016_ _0999_/X _1015_/X _1011_/B _1018_/B VSS VDD sky130_fd_sc_hd__or3_4
XANTENNA__1292__B1 _1254_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_262 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_34_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_295 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1595__A1 _1587_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1918_ _1843_/Y _1569_/B _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1849_ _1921_/D _1849_/LO VSS VDD sky130_fd_sc_hd__conb_1
XANTENNA__1595__B2 SCAN_IN[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_306 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_1_339 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1889__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1832__B _1828_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_207 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_44 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_346 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_229 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1807__C1 _1806_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_88 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1283__B1 _1254_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_417 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1279__B _1264_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_276 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_43_87 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1586__A1 _1120_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1338__A1 _1334_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_59 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1742__B _1695_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_73 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_0_350 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_48_365 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_398 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_63_357 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_232 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_3 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_290 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1703_ _1703_/A _1703_/B _1703_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1634_ _1597_/A _1633_/X _1597_/A _1633_/X _1634_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1329__A1 _1460_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1565_ _1812_/A _1769_/A _1575_/A _1564_/X _1566_/A VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_58_129 VSS VDD sky130_fd_sc_hd__fill_2
X_1496_ _1524_/B _1502_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_39_310 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_343 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_354 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1280__A3 _1259_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_287 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1827__B _1824_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_438 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1740__B2 _1739_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1740__A1 _1713_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_449 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_76 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_45_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_57_195 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_154 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_143 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_132 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1904__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_203 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1008__B1 _0977_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_74 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1737__B _1730_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1559__A1 _1905_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1559__B2 _1558_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_94 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1753__A _1753_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1350_ SCAN_IN[11] _1219_/X _1350_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1731__A1 _1729_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1472__B _1472_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1903__D _1740_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_180 VSS VDD sky130_fd_sc_hd__decap_6
X_1281_ _1279_/Y _1281_/B _1281_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_0_191 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_173 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_132 VSS VDD sky130_fd_sc_hd__decap_4
X_0996_ _0927_/X _1082_/D _0996_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_8_280 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1366__C _1366_/C VSS VDD sky130_fd_sc_hd__diode_2
X_1617_ _1616_/X _1617_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_5_91 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1663__A _1662_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1548_ _1619_/B _1548_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1722__A1 _1124_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_416 VSS VDD sky130_fd_sc_hd__decap_6
X_1479_ _1097_/X _1217_/A _1245_/A _1218_/A _1479_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1860__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_121 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1486__B1 _1475_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_324 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_357 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1838__A _1837_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_206 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_44 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1276__C _1276_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1573__A _1698_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_235 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1477__B1 _1476_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_121 VSS VDD sky130_fd_sc_hd__fill_1
X_1402_ _1897_/Q _1402_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_39_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_235 VSS VDD sky130_fd_sc_hd__decap_8
X_1333_ _1333_/A SCAN_IN[20] _1333_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_68_257 VSS VDD sky130_fd_sc_hd__decap_8
X_1264_ _1261_/Y _1263_/X _1261_/Y _1262_/Y _1264_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_452 VSS VDD sky130_fd_sc_hd__decap_6
X_1195_ _1897_/Q _1196_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_24_305 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1404__A2_N _1395_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_113 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_179 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1658__A _1546_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0994__A2 _0937_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1377__B _1376_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0979_ _1871_/Q _0932_/X _0933_/X _0979_/X VSS VDD sky130_fd_sc_hd__a21bo_4
XFILLER_10_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_25 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1393__A _1304_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_202 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_59_257 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1840__B _1837_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1474__A3 _1469_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_33 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_433 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_66 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1568__A _1630_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1631__B1 _1630_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_54 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1734__C _1716_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_9 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1750__B _1716_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_249 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_18_110 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_132 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_73_282 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_187 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1478__A _1417_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1622__B1 _1621_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1882_ _1450_/Y _1157_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
X_1316_ _1309_/X _1314_/X _1316_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1153__A2 _1149_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_419 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_227 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1660__B _1794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_249 VSS VDD sky130_fd_sc_hd__fill_2
X_1247_ _1247_/A _1525_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_260 VSS VDD sky130_fd_sc_hd__fill_2
X_1178_ _1461_/A _1167_/Y _1177_/X _1178_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_64_293 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_135 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_119 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_108 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_319 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1388__A _1241_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_341 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_374 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_13 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_46 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1835__B _1831_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1392__A2 _1386_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1144__A2 _1133_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1570__B _1705_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_282 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_422 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_433 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_252 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_620 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_53 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_631 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1604__B1 _1908_/Q VSS VDD sky130_fd_sc_hd__diode_2
XPHY_697 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_363 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_323 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_312 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_301 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1080__A1 _0964_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1080__B2 _0961_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0930__A _1868_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_367 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1745__B _1745_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_7 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1761__A _1763_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1135__A2 _1130_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1480__B _1334_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1911__D _1820_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1101_ _1097_/X _1245_/A _1100_/X _1101_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1032_ _0998_/A _1032_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_61_230 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1843__B1 _1502_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_296 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_127 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_149 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1001__A _0982_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1071__A1 _1871_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1865_ _1102_/Y _1865_/Q _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
X_1796_ _1181_/A _1796_/B _1796_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1374__A2 _1373_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_216 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1390__B _1390_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_282 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_252 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_466 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_436 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_8_109 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_160 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1846__A BB_IN VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_337 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1365__A2 _1364_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_149 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1581__A _1903_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_86 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_422 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_444 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_455 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0925__A _0925_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_425 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_450 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_7_131 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_120 VSS VDD sky130_fd_sc_hd__fill_2
X_1650_ _1575_/Y _1605_/X _1646_/Y _1649_/Y _1777_/C VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_11_193 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1906__D _1906_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1581_ _1903_/Q SCAN_IN[5] _1581_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1356__A2 _1351_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_171 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_293 VSS VDD sky130_fd_sc_hd__fill_2
X_1015_ _0968_/A _1015_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1292__A1 _1157_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1328__A1_N _1284_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1917_ _1839_/X _1567_/A _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1595__A2 SCAN_IN[2] VSS VDD sky130_fd_sc_hd__diode_2
X_1848_ _1713_/X _1813_/X _1064_/X _1848_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1779_ _1778_/A _1772_/X _1781_/B VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1878__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_300 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_67 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1807__B1 _1794_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1283__B2 _1282_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1283__A1 _1199_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_425 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1279__C _1278_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_469 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_266 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_288 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1576__A _1575_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1586__A2 _1265_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_145 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1338__A2 _1335_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_52 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_85 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_0_373 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_388 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_296 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_280 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_299 VSS VDD sky130_fd_sc_hd__fill_2
X_1702_ _1702_/A _1694_/B _1694_/C _1703_/B VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_69_3 VSS VDD sky130_fd_sc_hd__decap_6
X_1633_ _1729_/A _1263_/X _1596_/Y _1584_/X _1633_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1329__A2 _1326_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1564_ _1560_/X _1562_/X _1563_/X _1564_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1495_ _1492_/X _1524_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_39_300 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_322 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_174 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_358 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_62_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_299 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1856__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1396__A _1237_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1827__C _1825_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_148 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_428 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1740__A2 _1734_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1205__A1_N _1200_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_159 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_141 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_38_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_54_76 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1661__D1 _1660_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_277 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1008__A1 _1001_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_64 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1559__A2 _1557_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1753__B _1745_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1731__A2 _1719_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1192__B1 _1469_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1472__C _1472_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_439 VSS VDD sky130_fd_sc_hd__fill_2
X_1280_ _1127_/X SCAN_IN[4] _1259_/X _1259_/A SCAN_IN[5] _1281_/B VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_36_303 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_166 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_51_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_306 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1879__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_0995_ _0995_/A _0995_/B _0986_/X _0995_/D _1082_/D VSS VDD sky130_fd_sc_hd__nor4_4
XANTENNA__1366__D _1365_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1616_ _1594_/A _1615_/X _1594_/A _1615_/X _1616_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1634__A2_N _1633_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1547_ _1547_/A _1619_/B VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1722__A2 _1720_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1183__B1 _1182_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_428 VSS VDD sky130_fd_sc_hd__fill_2
X_1478_ _1417_/X _1349_/B _1478_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_74_409 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1486__A1 _1147_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_166 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_391 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_350 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1838__B _1836_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_424 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1477__A1 _1147_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_442 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_347 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1917__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_306 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_136 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_125 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_188 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1712__A1_N _1701_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_169 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_147 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__0933__A _1871_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1764__A _1763_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1401_ _1401_/A _1400_/Y _1401_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1914__D _1830_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_247 VSS VDD sky130_fd_sc_hd__decap_8
X_1332_ _1332_/A _1333_/A VSS VDD sky130_fd_sc_hd__inv_8
X_1263_ _1262_/Y _1263_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_431 VSS VDD sky130_fd_sc_hd__fill_1
X_1194_ _1113_/X _1188_/X _1193_/X _1194_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_36_144 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1004__A _0953_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_317 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_391 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_158 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_147 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_361 VSS VDD sky130_fd_sc_hd__fill_2
X_0978_ _0978_/A _0980_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1674__A _1674_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_48 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1393__B _1379_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_214 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_100 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_420 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_111 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_328 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_56 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_309 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_78 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1568__B _1544_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1631__A1 _1716_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_33 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0928__A _1874_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1750__C _1716_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_144 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_61_412 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1759__A _1759_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_158 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1478__B _1349_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1622__A1 _1546_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1909__D _1909_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1881_ _1441_/X _1146_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1917__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1494__A _1494_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1315_ _1309_/X _1314_/X _1216_/A _1315_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_56_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_93 VSS VDD sky130_fd_sc_hd__decap_3
X_1246_ _1240_/A _1247_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_49_280 VSS VDD sky130_fd_sc_hd__decap_4
X_1177_ _1463_/A _1166_/X _1177_/X VSS VDD sky130_fd_sc_hd__or2_4
XPHY_109 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_158 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1669__A SCAN_IN[14] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_331 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_386 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1392__A3 _1387_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_610 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1579__A _1579_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_643 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_632 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_106 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_687 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_76 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1604__A1 _1812_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1604__B2 _1286_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_698 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_375 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1080__A2 _1866_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_346 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0930__B _0929_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_353 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_331 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1761__B _1686_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1540__B1 _1539_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1100_ _1494_/A _1100_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_38_206 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_209 VSS VDD sky130_fd_sc_hd__decap_6
X_1031_ _1068_/B _1025_/X _1030_/X _1031_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_46_250 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_412 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1843__A1 _1652_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1071__A2 _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1864_ _1923_/Q _1065_/A _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1795_ _1089_/X _1658_/X _1795_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_29_206 VSS VDD sky130_fd_sc_hd__decap_4
X_1229_ _1228_/Y _1513_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_25_423 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1399__A _1398_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1598__B1 _1903_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_57 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_305 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_20_194 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_4_349 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_79_106 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1581__B SCAN_IN[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_76 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_356 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_31 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_231 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_404 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_415 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_253 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_448 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_440 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__A _0941_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_473 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VSS VDD sky130_fd_sc_hd__fill_2
X_1580_ _1741_/A _1256_/X _1741_/A _1256_/X _1580_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1772__A _1772_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_393 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1922__D _1922_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1014_ _1014_/A _1014_/B _1013_/X _1852_/D VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1292__A2 SCAN_IN[7] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1012__A _1011_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_459 VSS VDD sky130_fd_sc_hd__decap_8
X_1916_ _1916_/D _1609_/A _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1847_ _1847_/A _1847_/B _1847_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1595__A3 _1585_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1778_ _1778_/A _1751_/B _1778_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1854__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1482__A1_N _1103_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_378 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_356 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_24 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_72_337 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1807__A1 _1718_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1283__A2 _1579_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_404 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_253 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_234 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_256 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_301 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_153 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_164 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_337 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0936__A _0935_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_253 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_270 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_8_430 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1884__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_281 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1701_ _1587_/Y _1695_/B _1701_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1917__D _1839_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1632_ _1632_/A _1729_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1563_ _1186_/A _1796_/B _1181_/A _1608_/A _1563_/X VSS VDD sky130_fd_sc_hd__o22a_4
X_1494_ _1494_/A _1502_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_58_109 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1007__A _0980_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_337 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_54_326 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_315 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_304 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_197 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_392 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_429 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1827__D _1827_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1740__A3 _1735_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_56 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_164 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_189 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_329 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_54_44 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_201 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_223 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1587__A _1587_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_216 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1661__C1 _1659_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_21 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_289 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1008__A2 _1006_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1559__A3 _1539_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_98 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_411 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_444 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_79_63 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_68_407 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1192__A1 _1461_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1192__B2 _1177_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_451 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_178 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1497__A _1334_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0994_ _1061_/A _0937_/X _0991_/Y _0993_/X _0995_/D VSS VDD sky130_fd_sc_hd__a211o_4
X_1615_ _1587_/Y _1269_/Y _1614_/X _1615_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1546_ _1694_/A _1546_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_5_60 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1183__A1 _1771_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1477_ _1147_/A _1513_/A _1476_/X _1477_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_39_142 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_67_462 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1486__A2 _1513_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_189 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_215 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_362 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1200__A _1165_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_77 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1477__A2 _1513_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_337 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_98 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_65_87 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_156 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0933__B _0932_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_351 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1110__A _1110_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_230 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_53_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_285 VSS VDD sky130_fd_sc_hd__fill_2
X_1400_ _1304_/X _1397_/X _1399_/Y _1400_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1780__A _1778_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_215 VSS VDD sky130_fd_sc_hd__fill_2
X_1331_ _1525_/A _1288_/X _1468_/C _1382_/A VSS VDD sky130_fd_sc_hd__o21ai_4
X_1262_ SCAN_IN[4] _1262_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_64_410 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_76_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_443 VSS VDD sky130_fd_sc_hd__decap_3
X_1193_ _1833_/A _1193_/B _1193_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_36_178 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0979__A1 _1871_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_373 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1020__A _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_395 VSS VDD sky130_fd_sc_hd__fill_2
X_0977_ _0957_/Y _0970_/X _0972_/Y _0977_/D _0977_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1674__B _1661_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1529_ _1529_/A _1529_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1690__A _1690_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_237 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_292 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_67_281 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_432 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_402 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_13 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_104 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1568__C _1552_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_351 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1631__A2 _1616_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_255 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1869__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1105__A _1104_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_424 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0944__A _0951_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1759__B _1694_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_446 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_90 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1622__A2 _1590_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_384 VSS VDD sky130_fd_sc_hd__fill_2
X_1880_ _1880_/D _1259_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_41_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_192 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1648__A2_N _1647_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1925__D BB_IN VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_3 VSS VDD sky130_fd_sc_hd__decap_3
X_1314_ _1217_/A _1310_/Y _1274_/X _1313_/Y _1314_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_2_61 VSS VDD sky130_fd_sc_hd__decap_4
X_1245_ _1245_/A _1245_/B _1245_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1015__A _0968_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1176_ _1176_/A _1461_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_273 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1669__B _1805_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1074__B1 _1871_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1685__A _1690_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_398 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_443 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_56 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_243 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_11 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_611 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1579__B _1579_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_276 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_644 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_118 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_677 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_170 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_23_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1604__A2 SCAN_IN[10] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_699 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_343 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_28 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_358 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0939__A _0940_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1540__A1 _1161_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_432 VSS VDD sky130_fd_sc_hd__fill_2
X_1030_ _1013_/B _1029_/Y _0998_/A _1030_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_61_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1843__A2 _1837_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_118 VSS VDD sky130_fd_sc_hd__decap_4
X_1863_ _1113_/X _0925_/A _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1794_ _1108_/X _1794_/B _1794_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_69_376 VSS VDD sky130_fd_sc_hd__decap_12
X_1228_ _1198_/A _1228_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1295__B1 _1257_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_402 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_295 VSS VDD sky130_fd_sc_hd__fill_2
X_1159_ _1905_/Q _1579_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_52_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_107 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_12_129 VSS VDD sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_clk_0_0 clkbuf_0_clk_0_0/X _1853_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1598__A1 _1583_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1598__B2 SCAN_IN[5] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_140 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_14 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_317 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_79_118 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_75_346 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1665__A1_N _1364_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1907__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_240 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_402 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_251 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_54 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_243 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_430 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_166 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_7_144 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1772__B _1764_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_335 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_379 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_66_368 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_346 VSS VDD sky130_fd_sc_hd__decap_12
X_1013_ _0964_/A _1013_/B _1013_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1277__B1 _1114_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_265 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_427 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_438 VSS VDD sky130_fd_sc_hd__decap_4
X_1915_ _1833_/X _1567_/C _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_8_93 VSS VDD sky130_fd_sc_hd__decap_4
X_1846_ BB_IN _1846_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1777_ _1777_/A _1776_/Y _1777_/C _1777_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1894__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_151 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_69_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_324 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_36 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1807__A2 _1805_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1203__A _1202_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_221 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_298 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_409 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1440__B1 _1402_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_331 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_342 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_397 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_313 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1113__A _1100_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_265 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_382 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_287 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_260 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_271 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ _1529_/X _1694_/X _1695_/Y _1698_/Y _1699_/X _1899_/D VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_8_442 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1431__B1 _1412_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_90 VSS VDD sky130_fd_sc_hd__fill_2
X_1631_ _1716_/A _1616_/X _1630_/X _1631_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
X_1562_ _1812_/A _1796_/B _1181_/A _1608_/A _1562_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1493_ _1219_/X _1492_/X _1113_/X _1886_/D VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1007__B _0979_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1023__A _0955_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_202 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_257 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1670__B1 _1669_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1829_ _1798_/B _1824_/Y _1829_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_1_139 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1489__B1 _1176_/A VSS VDD sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_clk_0_16 clkbuf_0_clk_0_16/X _1887_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_57_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_57_176 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_316 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_349 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_168 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_235 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1661__B1 _1657_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_11 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_239 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1413__B1 _1412_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_75 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1108__A _1587_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1192__A2 _1167_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1309__A2_N _1270_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_349 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_198 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1778__A _1778_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_360 VSS VDD sky130_fd_sc_hd__decap_4
X_0993_ _0992_/X _0993_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1497__B _1218_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1404__B1 _1401_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1614_ _1614_/A _1589_/Y _1614_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1545_ _1552_/A _1794_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_5_50 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1183__A2 _1171_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_94 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1018__A _1014_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1476_ _1199_/A _1442_/A _1476_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_39_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_349 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_308 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1767__B1_N _1766_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1688__A _1688_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1643__B1 _1642_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_374 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_385 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_396 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_77_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_67 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_360 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1634__B1 _1597_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1295__A2_N _1281_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_264 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1233__A2_N _1332_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_91 VSS VDD sky130_fd_sc_hd__fill_1
X_1330_ _1247_/A _1288_/X _1326_/Y _1329_/Y _1468_/C VSS VDD sky130_fd_sc_hd__a211o_4
XANTENNA__1780__B _1772_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1261_ _1127_/A _1261_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1192_ _1461_/A _1167_/Y _1885_/Q _1469_/A _1177_/X _1193_/B VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_36_124 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_135 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_105 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_116 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1625__B1 _1702_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1801__A2_N _1734_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1301__A _1238_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0979__A2 _0932_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1020__B _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0976_ _0976_/A _0975_/X _0977_/D VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1674__C _1676_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_39 VSS VDD sky130_fd_sc_hd__fill_2
X_1528_ _1688_/A _1529_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_59_249 VSS VDD sky130_fd_sc_hd__decap_8
X_1459_ _1453_/Y _1458_/Y _1459_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_67_260 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_25 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_70_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_127 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1616__B1 _1594_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_138 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1211__A _1239_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1568__D _1694_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_76_65 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_124 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_241 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_105 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1759__C _1694_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_458 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_138 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1121__A _1120_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_341 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_374 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_80 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_91 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_396 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0960__A _1866_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1313_ _1217_/Y _1273_/X _1312_/X _1313_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_56_208 VSS VDD sky130_fd_sc_hd__fill_2
X_1244_ _1243_/X _1244_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_37_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_433 VSS VDD sky130_fd_sc_hd__fill_2
X_1175_ _1175_/A _1176_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_311 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1074__B2 _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1685__B _1689_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_38 VSS VDD sky130_fd_sc_hd__fill_2
X_0959_ _1865_/Q _0959_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1851__D _1851_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1206__A _1238_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_455 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_414 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_425 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_601 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_458 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_634 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_23 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_623 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_355 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_399 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0939__B _0940_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1116__A _1115_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1540__A2 _1638_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0955__A _0955_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_255 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1786__A _1620_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_288 VSS VDD sky130_fd_sc_hd__fill_2
X_1862_ _1063_/Y _0983_/A _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1867__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1793_ _1745_/A _1743_/A _1790_/X _1792_/Y _1803_/A VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_69_344 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1026__A _1014_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_388 VSS VDD sky130_fd_sc_hd__decap_12
X_1227_ _1147_/A _1361_/A _1213_/X _1226_/X _1227_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XFILLER_37_241 VSS VDD sky130_fd_sc_hd__decap_3
X_1158_ _1443_/A _1148_/Y _1157_/X _1158_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1295__B2 _1281_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1089_ _1091_/A _1089_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_40_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_119 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_428 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1696__A _1566_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1598__A2 SCAN_IN[4] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1859__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_185 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_4_329 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_75_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_314 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_57_67 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_73_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_66 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_266 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_428 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_420 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_163 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_123 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_497 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_81 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_384 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_185 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1277__A1 _1268_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1012_ _1011_/B _1013_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_19_263 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_74_391 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1277__B2 SCAN_IN[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_255 VSS VDD sky130_fd_sc_hd__fill_1
X_1914_ _1830_/X _1536_/A _1847_/X _1920_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1845_ _1777_/A _1842_/A _1502_/A _1844_/X _1820_/D _1845_/Y VSS VDD sky130_fd_sc_hd__a2111oi_4
X_1776_ _1683_/X _1776_/Y VSS VDD sky130_fd_sc_hd__inv_8
Xclkbuf_1_0__f_clk_0_16 clkbuf_0_clk_0_16/X _1886_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_16
XFILLER_57_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_328 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_200 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1863__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_233 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_461 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1440__A1 _1149_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_19 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_306 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_71_361 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_244 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_214 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_225 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_261 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_8_454 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1431__A1 _1429_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1630_ _1630_/A _1629_/X _1630_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1561_ _1567_/A _1608_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1492_ _1469_/A _1240_/A _1491_/X _1492_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1007__C _1007_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_314 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_347 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_358 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1304__A _1304_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_361 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1670__A1 SCAN_IN[19] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_247 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_28 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_269 VSS VDD sky130_fd_sc_hd__decap_6
X_1828_ _1798_/B _1824_/Y _1828_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1759_ _1759_/A _1694_/B _1694_/C _1762_/B VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_1_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1489__B2 _1460_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_47 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_clk_0_48_A clkbuf_0_clk_0_48/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1214__A _1214_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_339 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_72_147 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1661__A1 _1346_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_56 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1413__A1 _1410_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_79_87 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1192__A3 _1885_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_122 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_188 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_158 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0963__A _0963_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1778__B _1751_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1101__B1 _1100_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_394 VSS VDD sky130_fd_sc_hd__decap_3
X_0992_ _0992_/A _0990_/X _0992_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1404__B2 _1403_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1794__A _1108_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_291 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_3 VSS VDD sky130_fd_sc_hd__decap_4
X_1613_ _1613_/A _1805_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1168__B1 _1167_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1544_ _1544_/A _1613_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_5_62 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1018__B _1018_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1475_ _1157_/A _1516_/A _1138_/X _1361_/A _1475_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_280 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_111 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1034__A _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_328 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_158 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1643__A1 _1637_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_206 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_15 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1854__D _1022_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_438 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_46 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_12 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1331__B1 _1468_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0__f_clk_0_16_A clkbuf_0_clk_0_16/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_434 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_412 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_383 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1634__B2 _1633_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1119__A _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0958__A _1867_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1260_ _1430_/A _1258_/Y _1259_/X _1279_/A VSS VDD sky130_fd_sc_hd__o21ai_4
X_1191_ _1191_/A _1469_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_76_294 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_64_434 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1789__A _1789_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_158 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_17_361 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1625__A1 _1623_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1301__B _1299_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1020__C _1019_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1892__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_0975_ _1872_/Q _0933_/X _0934_/X _0975_/X VSS VDD sky130_fd_sc_hd__a21bo_4
XANTENNA__1389__B1 _1097_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1674__D _1673_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1029__A _1028_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_217 VSS VDD sky130_fd_sc_hd__fill_2
X_1527_ _1405_/X _1492_/X _1113_/X _1527_/X VSS VDD sky130_fd_sc_hd__o21a_4
X_1458_ _1421_/B _1456_/X _1457_/X _1458_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XANTENNA__1355__A2_N _1351_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_49 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1313__B1 _1312_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1389_ _1094_/X _1388_/X _1097_/X _1237_/A _1390_/B VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_70_415 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_37 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_48 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1616__B2 _1615_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_459 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_448 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1077__C1 _1061_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_250 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_423 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_158 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_73_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_404 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1402__A _1897_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_117 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_353 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_81 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_70 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_81 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_92 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_161 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1791__B1 _1161_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1312_ _1219_/A _1311_/X _1274_/A _1312_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_1243_ _1243_/A _1243_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_2_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_37_401 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_423 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_231 VSS VDD sky130_fd_sc_hd__fill_2
X_1174_ _1463_/A _1175_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_64_264 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_415 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_24_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_345 VSS VDD sky130_fd_sc_hd__fill_1
X_0958_ _1867_/Q _0958_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1888__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0975__B1_N _0934_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1782__B1 _1529_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_231 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_286 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_253 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_602 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_139 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_635 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_57 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_679 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_338 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1773__B1 _1727_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_9 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_401 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0955__B _0954_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_231 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_61_234 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1132__A _1131_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_61_245 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1786__B _1786_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1861_ _1861_/D _0940_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1792_ _1792_/A _1792_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1910__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1307__A _1307_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_367 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1026__B _1024_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1226_ _1138_/X _1212_/X _1225_/X _1226_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_52_201 VSS VDD sky130_fd_sc_hd__decap_12
X_1157_ _1157_/A _1147_/X _1157_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_37_275 VSS VDD sky130_fd_sc_hd__fill_1
X_1088_ _1064_/X _1066_/Y _1084_/X _1085_/X _1087_/Y _1851_/D VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1598__A3 _1581_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_131 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_49 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1862__D _1063_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1217__A _1217_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_220 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1873__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_34 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_426 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_448 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_212 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_43_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_459 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_410 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_421 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_131 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_454 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_60 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_93 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1127__A _1127_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_197 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_220 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_242 VSS VDD sky130_fd_sc_hd__fill_2
X_1011_ _0999_/X _1011_/B _1014_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1277__A2 SCAN_IN[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_297 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_223 VSS VDD sky130_fd_sc_hd__decap_3
X_1913_ _1913_/D _1630_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_8_84 VSS VDD sky130_fd_sc_hd__fill_2
X_1844_ _1575_/A _1844_/B _1844_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1775_ _1762_/A _1769_/Y _1770_/X _1773_/X _1774_/X _1907_/D VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1037__A _1013_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_164 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_27_16 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1264__A1_N _1261_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1209_ _1199_/A _1198_/X _1208_/X _1209_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_25_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_43_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1500__A _1216_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1857__D _1857_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1440__A2 _1388_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_355 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_0_377 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_381 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_71 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_251 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1410__A _1114_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_262 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_422 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_440 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_273 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_433 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1431__A2 _1430_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1560_ _1533_/X _1537_/X _1540_/Y _1556_/Y _1559_/Y _1560_/X VSS VDD sky130_fd_sc_hd__o41a_4
XFILLER_3_160 VSS VDD sky130_fd_sc_hd__fill_2
X_1491_ _1191_/A _1240_/A _1490_/X _1491_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_3_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_101 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_304 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_326 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1078__A2_N _1869_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_384 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_395 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1320__A _1320_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1670__A2 _1837_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_281 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_292 VSS VDD sky130_fd_sc_hd__fill_2
X_1827_ _1827_/A _1824_/Y _1825_/X _1827_/D _1913_/D VSS VDD sky130_fd_sc_hd__and4_4
X_1758_ _1713_/X _1750_/Y _1751_/X _1756_/X _1757_/X _1758_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
X_1689_ _1689_/A _1694_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_1_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_15 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_57_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_57_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_351 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_58 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_384 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_395 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1661__A2 _1569_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_259 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_281 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1413__A2 _1411_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_44 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_410 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_76_432 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1405__A _1384_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_112 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_307 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_48_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_63_104 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0963__B _0962_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1101__A1 _1097_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0991_ _0991_/A _0990_/X _0991_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_44_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_230 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1794__B _1794_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_252 VSS VDD sky130_fd_sc_hd__decap_8
X_1612_ _1790_/B _1611_/X _1612_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_8_296 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1168__A1 _1166_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1543_ _1736_/A _1543_/B _1543_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_5_41 VSS VDD sky130_fd_sc_hd__fill_2
X_1474_ _1402_/X _1468_/X _1469_/X _1472_/Y _1473_/X _1474_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1018__C _1017_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_410 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_79_292 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_67_432 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_123 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_39_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_167 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1034__B _1028_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1643__A2 _1641_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1050__A _1041_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_50_354 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_207 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_443 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1870__D _1153_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1331__A1 _1525_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_424 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_73_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_446 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_68 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_129 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_395 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_343 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_354 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_222 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_60 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_71 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_30_93 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_432 VSS VDD sky130_fd_sc_hd__decap_12
X_1190_ _1189_/Y _1191_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_76_262 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0974__A _0981_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1789__B _1786_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_351 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1625__A2 _1624_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_395 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_365 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1020__D _1011_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_398 VSS VDD sky130_fd_sc_hd__fill_2
X_0974_ _0981_/A _0976_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1389__B2 _1237_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1389__A1 _1094_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1616__A1_N _1594_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1010__B1 _1061_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1526_ _1525_/A _1524_/C _1525_/Y _1064_/X _1492_/X _1896_/D VSS VDD sky130_fd_sc_hd__a2111oi_4
XANTENNA__1045__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_17 VSS VDD sky130_fd_sc_hd__fill_2
X_1457_ _1168_/X _1388_/X _1897_/Q _1457_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1313__A1 _1217_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1388_ _1241_/A _1388_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_55_424 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_104 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_148 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_70_405 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1077__B1 _0940_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_170 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_343 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_365 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_23_376 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1865__D _1102_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_56 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_262 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_435 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_61_416 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_438 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_60 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_71 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_82 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_151 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_184 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_195 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1791__A1 _1745_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1791__B2 _1790_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1311_ _1271_/A SCAN_IN[0] _1311_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1242_ _1245_/A _1245_/B _1243_/A VSS VDD sky130_fd_sc_hd__or2_4
X_1173_ _1827_/A _1168_/X _1107_/X _1172_/X _1173_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_49_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_195 VSS VDD sky130_fd_sc_hd__fill_1
X_0957_ _0957_/A _0957_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1231__B1 _1230_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1782__A1 _1188_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1857__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1509_ _1506_/X _1502_/B _1507_/Y _1509_/D _1890_/D VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__1298__B1 _1278_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1503__A _1307_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_257 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_625 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_306 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1222__B1 _1220_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1773__A1 _1771_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_78_335 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_413 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1882__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_446 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_243 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_46_254 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_276 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1132__B _1123_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_427 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_287 VSS VDD sky130_fd_sc_hd__decap_12
X_1860_ _1860_/D _1860_/Q _1847_/X _1865_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1791_ _1745_/A _1743_/A _1161_/A _1790_/B _1792_/A VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_42_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_324 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1307__B _1306_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1026__C _1025_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_221 VSS VDD sky130_fd_sc_hd__fill_2
X_1225_ _1127_/X _1307_/A _1222_/X _1224_/X _1225_/X VSS VDD sky130_fd_sc_hd__o22a_4
X_1156_ _1199_/A _1443_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_52_213 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_52_257 VSS VDD sky130_fd_sc_hd__fill_2
X_1087_ _1085_/A CLK_OUT _1833_/A _1087_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_20_154 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1906__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_46 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_276 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_400 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_408 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_411 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_290 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_110 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_455 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_143 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_7_114 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_488 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_176 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1746__A1 _1745_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_169 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1408__A _1342_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_397 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_305 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1143__A _1736_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1010_ _0985_/A _0942_/A _1009_/X _1061_/A _0937_/X _1011_/B VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_47_91 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1277__A3 _1266_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1682__B1 _1673_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1293__A2_N _1292_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_290 VSS VDD sky130_fd_sc_hd__fill_1
X_1912_ _1823_/Y _1544_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_30_441 VSS VDD sky130_fd_sc_hd__fill_2
X_1843_ _1652_/Y _1837_/X _1502_/A _1844_/B _1820_/D _1843_/Y VSS VDD sky130_fd_sc_hd__a2111oi_4
X_1774_ _1183_/X _1709_/A _1529_/A _1774_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1318__A _1307_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1037__B _1082_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_143 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_69_176 VSS VDD sky130_fd_sc_hd__decap_3
X_1208_ _1166_/A _1516_/A _1208_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1053__A _0940_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1139_ _1138_/X _1128_/X _1139_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_13_408 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_419 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1425__B1 _1196_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_238 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1500__B _1498_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_106 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1873__D _1184_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1228__A _1198_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_367 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_389 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_327 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_75_168 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_75_157 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_83 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1920__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_396 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_252 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1410__B _1399_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_263 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_82 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_8_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1138__A _1259_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1490_ _1461_/A _1460_/A _1488_/X _1489_/X _1490_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__0977__A _0957_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_168 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_54_319 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_308 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1655__B1 SCAN_IN[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_205 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1320__B _1300_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_290 VSS VDD sky130_fd_sc_hd__decap_3
X_1826_ _1813_/X _1827_/D VSS VDD sky130_fd_sc_hd__inv_8
X_1757_ _1163_/X _1709_/A _1529_/A _1757_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1048__A _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1688_ _1688_/A _1703_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_38_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_72_105 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_48 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1511__A _1361_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1868__D _1135_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_56 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_82 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_179 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_138 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1637__B1 _1636_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_393 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_341 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1421__A _1130_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1101__A2 _1245_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_71_171 VSS VDD sky130_fd_sc_hd__fill_1
X_0990_ _1873_/Q _0934_/X _0936_/Y _0990_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_12_260 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_80 VSS VDD sky130_fd_sc_hd__decap_12
X_1611_ _1600_/X _1610_/X _1600_/X _1610_/X _1611_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1168__A2 _1157_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1542_ _1630_/A _1543_/B VSS VDD sky130_fd_sc_hd__inv_8
X_1473_ _1193_/B _1401_/A _1196_/A _1473_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_67_400 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_39_135 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_352 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1050__B _1045_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_311 VSS VDD sky130_fd_sc_hd__decap_8
X_1809_ _1803_/A _1808_/Y _1792_/A _1790_/X _1809_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1506__A _1100_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_433 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_455 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1331__A2 _1288_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_308 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_65_36 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_352 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1241__A _1241_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_322 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_377 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_73 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_5_245 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_5_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_267 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_219 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1416__A _1349_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_444 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_76_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_274 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1789__C _1787_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_330 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_190 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_127 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1151__A _1150_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_182 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_377 VSS VDD sky130_fd_sc_hd__fill_2
X_0973_ _0973_/A _0981_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1389__A2 _1388_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1010__B2 _0937_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1010__A1 _0985_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1525_ _1525_/A _1524_/C _1525_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1326__A _1460_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1045__B _1044_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1456_ _1452_/A _1447_/A _1463_/B _1456_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_67_230 VSS VDD sky130_fd_sc_hd__decap_8
X_1387_ _1097_/X _1379_/B _1387_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XFILLER_67_285 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1313__A2 _1273_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_447 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1061__A _1061_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1077__A1 _0973_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_160 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_119 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_355 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_196 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1881__D _1441_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_259 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_58_241 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_58_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_46_414 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_73_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_266 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_61_428 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_322 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_50 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_61 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_72 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_83 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_388 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_94 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_94 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1791__A2 _1743_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_8 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1146__A _1146_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1310_ _1273_/X _1310_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_1_270 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0985__A _0985_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_43 VSS VDD sky130_fd_sc_hd__fill_2
X_1241_ _1241_/A _1397_/C _1245_/B VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1584__A2_N _1263_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1172_ _1169_/X _1162_/X _1171_/Y _1172_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_2_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_255 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_24_108 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_60_450 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_163 VSS VDD sky130_fd_sc_hd__decap_12
X_0956_ _0955_/X _0957_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1231__A1 _1199_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1782__A2 _1709_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1537__A2_N _1609_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0990__B1 _0936_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1056__A _1058_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1508_ _1212_/X _1503_/X _1509_/D VSS VDD sky130_fd_sc_hd__or2_4
X_1439_ _1401_/A _1438_/Y _1439_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1897__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1298__A1 _1261_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_222 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_425 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1298__B2 _1264_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1503__B _1501_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_428 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_247 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_626 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_303 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1876__D _1392_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_347 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_196 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_329 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1222__B2 _1221_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1222__A1 _1114_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1773__A2 _1772_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_74 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_211 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_46_266 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_439 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_60 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_299 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_130 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_174 VSS VDD sky130_fd_sc_hd__decap_12
X_1790_ _1753_/A _1790_/B _1790_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_52_81 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_69_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_358 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_69_347 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_391 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_37_233 VSS VDD sky130_fd_sc_hd__decap_8
X_1224_ _1115_/Y _1394_/A _1127_/X _1215_/A _1224_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1155_ _1155_/A _1199_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_25_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_255 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_19 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_439 VSS VDD sky130_fd_sc_hd__fill_2
X_1086_ _1923_/Q _1833_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_37_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_144 VSS VDD sky130_fd_sc_hd__fill_2
X_0939_ _0940_/A _0940_/B _0995_/A VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_75_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1514__A _1513_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_380 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_266 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1140__B1 _1139_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_401 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_450 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_412 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_269 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_1_0_A _CTS_root/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_445 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_155 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_478 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_148 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1746__A2 _1745_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_343 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1408__B _1408_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_111 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_177 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_317 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_9 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1143__B _1132_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_277 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1682__A1 _1675_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_34_247 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_258 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_91 VSS VDD sky130_fd_sc_hd__fill_2
X_1911_ _1820_/Y _1552_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_30_420 VSS VDD sky130_fd_sc_hd__decap_3
X_1842_ _1842_/A _1844_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_8_53 VSS VDD sky130_fd_sc_hd__decap_8
X_1773_ _1771_/X _1772_/X _1727_/X _1773_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_8_97 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1318__B _1308_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1370__B1 _1338_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1334__A _1217_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_309 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_65_350 VSS VDD sky130_fd_sc_hd__fill_2
X_1207_ _1352_/A _1516_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_372 VSS VDD sky130_fd_sc_hd__decap_12
X_1138_ _1259_/A _1138_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1069_ _1872_/Q _1040_/X _1067_/X _1068_/X _1082_/A VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_25_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_206 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_28 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1425__A1 _1421_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1872__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1509__A _1506_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_302 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_68_58 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_36 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_75_103 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1244__A _1243_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__CTS_buf_1_0_A _CTS_buf_1_0/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_361 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_203 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_394 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_353 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_95 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_31_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_386 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_242 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_413 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_264 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_297 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_94 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1419__A _1417_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1306__A2_N _1305_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0927__B1 _1065_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_184 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0977__B _0970_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1154__A _1157_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0993__A _0992_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_350 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1655__B2 _1558_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_375 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1320__C _1319_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_239 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1895__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_1825_ _1724_/A _1822_/X _1825_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1756_ _1752_/X _1755_/Y _1727_/X _1756_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1048__B _1037_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1687_ _1571_/A _1695_/B _1687_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1064__A _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1343__B1 _1394_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_372 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_364 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1511__B _1509_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1884__D _1466_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1239__A _1239_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1582__B1 _1581_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_187 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1702__A _1702_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1637__A1 _1627_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1421__B _1421_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_71 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_93 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1610_ _1905_/Q SCAN_IN[7] _1579_/X _1610_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_8_276 VSS VDD sky130_fd_sc_hd__fill_2
X_1541_ _1536_/A _1798_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_5_54 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0988__A _1860_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_98 VSS VDD sky130_fd_sc_hd__fill_2
X_1472_ _1412_/X _1472_/B _1472_/C _1472_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_79_261 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_67_423 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1612__A _1790_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_117 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1813__A2_N _1812_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_191 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_150 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_183 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_389 VSS VDD sky130_fd_sc_hd__fill_1
X_1808_ _1804_/Y _1805_/X _1807_/X _1800_/A _1801_/X _1808_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
XANTENNA__1059__A _1032_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1739_ _1144_/X _1720_/X _1529_/X _1739_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1564__B1 _1563_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1910__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_38 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_65_48 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1522__A _1333_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_117 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_331 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1879__D _1879_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_364 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1241__B _1397_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_334 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_367 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_52 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_85 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1555__B1 _1554_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_257 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1879__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1416__B _1408_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_423 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1789__D _1788_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_448 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_320 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_70 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_51_109 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_312 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_334 VSS VDD sky130_fd_sc_hd__fill_2
X_0972_ _0971_/Y _0972_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_32_389 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_91 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_65_3 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1607__A _1601_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1010__A2 _0942_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1524_ _1100_/X _1524_/B _1524_/C _1524_/D _1895_/D VSS VDD sky130_fd_sc_hd__and4_4
XANTENNA__1326__B _1326_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1455_ _1462_/B _1463_/B VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_67_242 VSS VDD sky130_fd_sc_hd__fill_2
X_1386_ _1334_/X _1383_/B _1386_/C _1386_/X VSS VDD sky130_fd_sc_hd__or3_4
XFILLER_55_415 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1342__A _1342_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1061__B _1061_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_109 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_429 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1077__A2 _1076_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_323 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_367 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_39 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1537__B1 _1741_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1517__A _1516_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_58_220 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_212 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1252__A _1200_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_73_245 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_109 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_40 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_62 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_51 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_62 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_73 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_378 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_73 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_84 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_95 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_83 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1427__A _1427_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_282 VSS VDD sky130_fd_sc_hd__fill_2
X_1240_ _1240_/A _1240_/B _1240_/C _1239_/X _1397_/C VSS VDD sky130_fd_sc_hd__nor4_4
XFILLER_49_242 VSS VDD sky130_fd_sc_hd__fill_2
X_1171_ _1170_/X _1171_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_37_415 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1700__B1 _1698_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1162__A _1905_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_99 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_37_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_407 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_418 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_175 VSS VDD sky130_fd_sc_hd__decap_12
X_0955_ _0955_/A _0954_/Y _0955_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1231__A2 _1205_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_382 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0990__A1 _1873_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1337__A SCAN_IN[11] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1056__B _1060_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1507_ _1212_/X _1503_/X _1507_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1438_ _1434_/A _1430_/X _1437_/X _1438_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XANTENNA__1298__A2 _1263_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1369_ _1369_/A _1369_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_55_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_70_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1800__A _1800_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_418 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_616 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_605 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_649 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_49 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_38 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_627 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_315 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1758__B1 _1756_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1222__A2 _1216_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1892__D _1515_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_53 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1247__A _1247_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_86 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_78_337 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_46_223 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1710__A _1688_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_186 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_93 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1749__B1 _1747_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_381 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_363 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1157__A _1157_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_315 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0996__A _0927_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_3 VSS VDD sky130_fd_sc_hd__decap_3
X_1223_ _1216_/A _1394_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1154_ _1157_/A _1155_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_37_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_215 VSS VDD sky130_fd_sc_hd__fill_2
X_1085_ _1085_/A _1084_/B _1085_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_37_278 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1620__A _1092_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0938_ _0928_/Y _0936_/Y _0937_/X _0940_/B VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1067__A _1023_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_318 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_57_27 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1514__B _1511_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_392 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1140__A1 _1430_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_15 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_429 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1530__A _1569_/B VSS VDD sky130_fd_sc_hd__diode_2
XPHY_402 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1887__D _1499_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_123 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_446 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_479 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_52 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_85 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0954__A1 _1868_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1408__C _1408_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_355 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1705__A _1093_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_189 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_329 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_289 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_215 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_395 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1682__A2 _1681_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_462 VSS VDD sky130_fd_sc_hd__decap_8
X_1910_ _1910_/D _1694_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_42_270 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_8_32 VSS VDD sky130_fd_sc_hd__decap_6
X_1841_ _1840_/X _1842_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1772_ _1772_/A _1764_/Y _1772_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__0945__A1 _1869_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1318__C _1317_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_156 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1370__A1 _1334_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1206_ _1238_/B _1352_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_65_384 VSS VDD sky130_fd_sc_hd__decap_12
X_1137_ _1259_/A _1430_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_25_204 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1350__A SCAN_IN[11] VSS VDD sky130_fd_sc_hd__diode_2
X_1068_ _1870_/Q _1068_/B _1068_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1425__A2 _1424_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1509__B _1502_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_26 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1525__A _1525_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1629__A1_N _1596_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_373 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_332 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_210 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_410 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_243 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_254 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1419__B _1419_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0927__B2 _1494_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_196 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1435__A _1198_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0977__C _0972_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_126 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_318 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_329 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1170__A _1169_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1475__A2_N _1516_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_384 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_91 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_62_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_240 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_30_262 VSS VDD sky130_fd_sc_hd__fill_2
X_1824_ _1724_/A _1822_/X _1824_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1755_ _1754_/X _1755_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1686_ _1686_/A _1695_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1343__A1 _1342_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1343__B2 _1339_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_137 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_376 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_428 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_417 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1239__B _1214_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1031__B1 _1030_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1582__A1 _1737_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1255__A SCAN_IN[6] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1553__A1_N _1120_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_402 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_104 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_126 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_76_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1702__B _1694_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1637__A2 _1631_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_310 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_162 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_398 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_83 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1270__B1 _1304_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_288 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_93 VSS VDD sky130_fd_sc_hd__fill_2
X_1540_ _1161_/A _1638_/A _1539_/X _1540_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_5_22 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_450 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1165__A _1165_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1471_ _1469_/A _1471_/B _1472_/C VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_79_273 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1325__A1 _1451_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_104 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_115 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_3 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1612__B _1611_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1862__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_321 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_346 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1797__D1 _1796_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1807_ _1718_/A _1805_/B _1794_/X _1806_/X _1807_/X VSS VDD sky130_fd_sc_hd__a211o_4
XANTENNA__1059__B _1057_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1738_ _1736_/X _1745_/B _1720_/X _1738_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1564__A1 _1560_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1075__A _1071_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1669_ SCAN_IN[14] _1805_/B _1669_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_49_28 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1803__A _1803_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_416 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_73_449 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_438 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1522__B _1523_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_398 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1895__D _1895_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1555__A1 _1736_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_85 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_420 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1416__C _1408_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1713__A _1703_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1885__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_72 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_276 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_64_427 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_170 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_82 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_17_365 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_387 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_151 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1491__B1 _1490_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0971_ _0955_/A _0954_/Y _0963_/A _0962_/X _0971_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XANTENNA__0999__A _0964_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1913__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1607__B _1607_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1010__A3 _1009_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1523_ _1333_/A _1523_/B _1524_/D VSS VDD sky130_fd_sc_hd__nand2_4
X_1454_ _1452_/A _1447_/A _1462_/B VSS VDD sky130_fd_sc_hd__or2_4
X_1385_ _1196_/X _1244_/Y _1245_/X _1379_/X _1384_/X _1875_/D VSS VDD sky130_fd_sc_hd__o32ai_4
XFILLER_27_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1342__B _1341_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_184 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1482__B1 _1116_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1885__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_50_165 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1234__B1 _1176_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1537__B2 _1734_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_206 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_228 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1517__B _1516_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_232 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_58_210 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1533__A _1161_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_276 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1252__B _1578_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_302 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_30 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_41 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1473__B1 _1196_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_52 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_195 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_63 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_74 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_110 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_85 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_165 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_85 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_96 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1225__B1 _1222_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1427__B _1408_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1443__A _1443_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_23 VSS VDD sky130_fd_sc_hd__fill_1
X_1170_ _1169_/X _1162_/X _1170_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_2_67 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1700__A1 _1529_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1700__B2 _1699_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_70 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1162__B _1150_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_235 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_151 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1464__B1 _1421_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1900__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_187 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_198 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1767__A1 _1727_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0954_ _1868_/Q _0929_/X _0930_/X _0954_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XANTENNA__1231__A3 _1209_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1618__A _1590_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0990__A2 _0934_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1337__B _1219_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1506_ _1100_/X _1506_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1437_ _1434_/A _1430_/X _1437_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1353__A _1352_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1368_ _1366_/A _1368_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_46_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_257 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_235 VSS VDD sky130_fd_sc_hd__decap_4
X_1299_ _1279_/A _1298_/X _1279_/A _1298_/X _1299_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XPHY_617 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_606 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1758__A1 _1713_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1758__B2 _1757_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1528__A _1688_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_98 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_78_349 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_405 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1263__A _1262_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_449 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_216 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1923__CLK _1923_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_238 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_36_84 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_441 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1749__B2 _1748_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1157__B _1147_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_386 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0996__B _1082_/D VSS VDD sky130_fd_sc_hd__diode_2
X_1222_ _1114_/X _1216_/Y _1220_/X _1221_/X _1222_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_77_371 VSS VDD sky130_fd_sc_hd__fill_2
X_1153_ _1827_/A _1149_/X _1107_/X _1152_/X _1153_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_25_419 VSS VDD sky130_fd_sc_hd__fill_2
X_1084_ _1084_/A _1084_/B _1084_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1620__B _1619_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_290 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_441 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_135 VSS VDD sky130_fd_sc_hd__decap_3
X_0937_ _1874_/Q _0935_/X _0937_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1348__A _1239_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1067__B _1869_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1083__A CLK_OUT VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_202 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_73_27 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1140__A2 _1129_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_216 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_227 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_403 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_282 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_271 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_436 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_168 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_139 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1258__A SCAN_IN[5] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1600__B1 _1580_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_75 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_301 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0954__A2 _0929_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_78_135 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1705__B _1705_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_382 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_360 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_74_330 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1667__B1 _1346_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_83 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_290 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_11 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_30_433 VSS VDD sky130_fd_sc_hd__fill_2
X_1840_ _1652_/Y _1837_/X _1840_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1771_ _1771_/A _1763_/X _1771_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_8_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0945__A2 _0930_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1370__A2 _1335_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1205_ _1200_/Y _1442_/A _1434_/A _1427_/A _1205_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1136_ _1100_/X _1820_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_396 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_25_216 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_249 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1350__B _1219_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1067_ _1023_/Y _1869_/Q _1067_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_33_282 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1509__C _1507_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_315 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1525__B _1524_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_319 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1541__A _1536_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1898__D _1898_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_53 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_200 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_75 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_233 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_422 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_255 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_41 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_288 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_3_120 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1716__A _1716_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_164 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1435__B _1383_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0977__D _0977_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_466 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_60 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_330 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1451__A _1451_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1170__B _1162_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_388 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_252 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_296 VSS VDD sky130_fd_sc_hd__decap_4
X_1823_ _1820_/A _1821_/Y _1822_/X _1820_/D _1823_/Y VSS VDD sky130_fd_sc_hd__nor4_4
X_1754_ _1754_/A _1754_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1685_ _1690_/A _1689_/A _1686_/A VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1626__A _1623_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_105 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1343__A2 _1341_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_149 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1361__A _1361_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_341 VSS VDD sky130_fd_sc_hd__decap_4
X_1119_ _1923_/Q _1119_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_13_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_17 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_252 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_285 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1239__C _1216_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_15 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1031__A1 _1068_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1582__A2 _1258_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1536__A _1536_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_156 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_108 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1271__A _1271_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_63 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_341 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_363 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1702__C _1694_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_344 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_40 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_44_377 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_71_196 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_263 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_252 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1270__B2 _1269_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_223 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_61 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_267 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1446__A _1445_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_67 VSS VDD sky130_fd_sc_hd__decap_12
X_1470_ _1469_/A _1471_/B _1472_/B VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_69_92 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1325__A2 _1291_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_436 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_138 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_149 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1181__A _1181_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_333 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1797__C1 _1795_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1806_ _1795_/X _1787_/X _1788_/X _1806_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1059__C _1058_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1737_ _1737_/A _1730_/A _1745_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1564__A2 _1562_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1668_ _1567_/A _1837_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1075__B _1072_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1599_ _1597_/Y _1598_/X _1599_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1803__B _1797_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_447 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1091__A _1091_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_428 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_141 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_174 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_358 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_237 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1266__A _1114_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1555__A2 _1543_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_40 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_211 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1489__A2_N _1359_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_458 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_266 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_50 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_182 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1491__A1 _1191_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_369 VSS VDD sky130_fd_sc_hd__fill_2
X_0970_ _0964_/A _1865_/Q _0963_/Y _0969_/X _0970_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_71_71 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1176__A _1176_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1522_ _1333_/A _1523_/B _1524_/C VSS VDD sky130_fd_sc_hd__or2_4
X_1453_ _1402_/X _1451_/Y _1453_/C _1453_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_4_281 VSS VDD sky130_fd_sc_hd__decap_12
X_1384_ _1384_/A _1384_/B _1384_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_67_266 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_277 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_70_409 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_347 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1482__B2 _1342_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1234__B2 _1451_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1234__A1 _1189_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_177 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1086__A _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_16 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1533__B _1638_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_299 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_450 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_20 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_31 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_20 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_26_163 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_42 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1473__A1 _1193_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_53 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_53 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_64 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_75 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_86 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_97 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1225__B2 _1224_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1225__A1 _1127_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_188 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1852__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1427__C _1408_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1724__A _1724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_13 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_200 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1443__B _1419_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_255 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1700__A2 _1694_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_203 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_37_428 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_49_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_93 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_64_269 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1464__A1 _1462_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_122 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_32_144 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1767__A2 _1765_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_340 VSS VDD sky130_fd_sc_hd__fill_2
X_0953_ _1068_/B _0945_/X _1005_/A _0952_/Y _0953_/X VSS VDD sky130_fd_sc_hd__a211o_4
XFILLER_70_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1231__A4 _1227_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1505_ _1502_/A _1502_/B _1503_/X _1504_/Y _1505_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1436_ _1384_/A _1436_/B _1436_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1367_ _1338_/X _1345_/X _1357_/X _1366_/Y _1367_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1152__B1 _1151_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_439 VSS VDD sky130_fd_sc_hd__fill_2
X_1298_ _1261_/Y _1263_/X _1278_/Y _1264_/X _1298_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_70_228 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_607 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_420 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_62_29 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_629 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_188 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1758__A2 _1750_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1875__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0966__B1 _0961_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1875__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_11 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_44 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1544__A _1544_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1391__B1 _1384_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1901__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_203 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_54_280 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_431 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1719__A _1719_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_73 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_306 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1454__A _1452_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_81 VSS VDD sky130_fd_sc_hd__fill_1
X_1221_ _1103_/X _1217_/Y _1221_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_77_361 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1134__B1 _1133_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_203 VSS VDD sky130_fd_sc_hd__fill_1
X_1152_ _1904_/Q _1143_/X _1151_/Y _1152_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_37_225 VSS VDD sky130_fd_sc_hd__fill_2
X_1083_ CLK_OUT _1082_/Y _1084_/B VSS VDD sky130_fd_sc_hd__xnor2_4
XFILLER_37_269 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_52_239 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1898__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_272 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_114 VSS VDD sky130_fd_sc_hd__fill_2
X_0936_ _0935_/X _0936_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_9_192 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1373__B1 _1355_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1364__A SCAN_IN[16] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1083__B _1082_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1419_ _1417_/X _1419_/B _1419_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_68_372 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1125__B1 _1119_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_236 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_420 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_404 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_294 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_32 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1539__A _1169_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1600__A1 _1741_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1600__B2 _1599_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1274__A _1274_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_78_125 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_236 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1667__B2 _1569_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1667__A1 _1675_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_375 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_95 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_228 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_250 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_445 VSS VDD sky130_fd_sc_hd__decap_12
X_1770_ _1771_/A _1751_/B _1770_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_30_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_195 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_103 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1355__B1 _1352_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_147 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_180 VSS VDD sky130_fd_sc_hd__decap_3
X_1204_ _1238_/D _1427_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1135_ _1827_/A _1130_/X _1107_/X _1728_/A _1135_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_25_239 VSS VDD sky130_fd_sc_hd__fill_1
X_1066_ _1084_/A CLK_OUT _1066_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_21_445 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1359__A _1359_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1899_ _1899_/D _1091_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1509__D _1509_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1913__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1094__A _1094_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1822__A _1544_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_320 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1649__A1 _1769_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_386 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_367 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_201 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_234 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_445 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_267 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1890__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1269__A SCAN_IN[2] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_467 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_278 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_438 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1716__B _1716_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_143 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_412 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1435__C _1386_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_180 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1451__B _1383_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_323 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_312 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_74_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1179__A _1772_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1822_ _1544_/A _1821_/B _1822_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1753_ _1753_/A _1745_/X _1754_/A VSS VDD sky130_fd_sc_hd__or2_4
X_1684_ SCAN_IN[21] _1777_/A _1683_/X _1689_/A VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1626__B _1624_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1328__B1 _1284_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_117 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0927__A2_N _1494_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_128 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_320 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1361__B SCAN_IN[16] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_19 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_301 VSS VDD sky130_fd_sc_hd__decap_4
X_1118_ _1116_/X _1105_/Y _1117_/X _1118_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_53_367 VSS VDD sky130_fd_sc_hd__fill_2
X_1049_ _1032_/X _1047_/Y _1048_/X _1859_/D VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_0_90 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1089__A _1091_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_264 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1868__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1239__D _1217_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_27 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1031__A2 _1025_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_426 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_168 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1552__A _1552_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1271__B SCAN_IN[0] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_375 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_397 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1074__A2_N _1867_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_356 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_389 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_63 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_231 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_51 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1727__A _1696_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_79 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_69_60 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_67_415 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1462__A _1461_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_62_142 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_164 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_35_367 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_186 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_337 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1797__B1 _1794_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1805_ _1718_/A _1805_/B _1805_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1736_ _1736_/A _1730_/Y _1736_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1549__B1 _1089_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1667_ _1675_/A _1608_/A _1346_/Y _1569_/B _1673_/A VSS VDD sky130_fd_sc_hd__o22a_4
X_1598_ _1583_/A SCAN_IN[4] _1581_/X _1903_/Q SCAN_IN[5] _1598_/X VSS VDD sky130_fd_sc_hd__a32o_4
XANTENNA__1075__C _1073_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1721__B1 _1720_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1803__C _1803_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_437 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_109 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_164 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_11 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_41_326 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1788__B1 _1108_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_55 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1547__A _1547_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_21 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_32 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1266__B SCAN_IN[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_54 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1438__B1_N _1437_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_404 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1712__B1 _1709_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_52 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_194 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_131 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_367 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_164 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1491__A2 _1240_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_186 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_381 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_72_7 VSS VDD sky130_fd_sc_hd__decap_8
X_1521_ _1506_/X _1524_/B _1521_/C _1523_/B _1521_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1452_ _1452_/A _1378_/A _1453_/C VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_4_293 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_201 VSS VDD sky130_fd_sc_hd__fill_2
X_1383_ _1218_/A _1383_/B _1386_/C _1384_/B VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_67_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_407 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1922__RESET_B RESET_N VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_440 VSS VDD sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clk_1_0 clkbuf_0_clk_1_0/X _CTS_buf_1_32/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_63_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_315 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_175 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_359 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1234__A2 _1332_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_381 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1367__A _1338_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1719_ _1719_/A _1706_/X _1719_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_76_39 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_28 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_73_237 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1830__A _1827_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_21 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_10 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_315 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_337 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_32 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_43 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1473__A2 _1401_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_54 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_65 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_123 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_76 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_87 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_98 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1225__A2 _1307_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_381 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1724__B _1716_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_223 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1700__A3 _1695_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_131 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_440 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_281 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1464__A2 _1471_/B VSS VDD sky130_fd_sc_hd__diode_2
X_0952_ _0950_/X _0947_/X _0951_/X _0952_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1187__A _1812_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0975__A1 _1872_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1504_ _1307_/A _1501_/X _1504_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1435_ _1198_/X _1383_/B _1386_/C _1436_/B VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1152__A1 _1904_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1366_ _1366_/A _1361_/X _1366_/C _1365_/X _1366_/Y VSS VDD sky130_fd_sc_hd__nand4_4
XFILLER_28_407 VSS VDD sky130_fd_sc_hd__decap_12
X_1297_ _1228_/Y _1297_/B _1320_/A VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_70_207 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_608 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_145 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1758__A3 _1751_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0966__A1 _1865_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1097__A _1096_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1825__A _1724_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_307 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1391__A1 _1243_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_134 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_52 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1719__B _1706_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_362 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_333 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_322 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1735__A _1737_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1454__B _1447_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_7 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_71 VSS VDD sky130_fd_sc_hd__fill_2
X_1220_ _1103_/X _1217_/Y _1094_/X _1219_/X _1220_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1134__A1 _1131_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1151_ _1150_/X _1151_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1470__A _1469_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1082_ _1082_/A _1075_/X _1081_/X _1082_/D _1082_/Y VSS VDD sky130_fd_sc_hd__nor4_4
XFILLER_20_148 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_160 VSS VDD sky130_fd_sc_hd__fill_2
X_0935_ _1873_/Q _0934_/X _0935_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1373__A1 _1369_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1373__B2 _1354_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_19 VSS VDD sky130_fd_sc_hd__fill_2
X_1418_ _1378_/A _1419_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1125__B2 _1124_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1125__A1 _1113_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1380__A _1897_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_215 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_248 VSS VDD sky130_fd_sc_hd__fill_1
X_1349_ _1347_/Y _1349_/B _1349_/X VSS VDD sky130_fd_sc_hd__and2_4
XPHY_405 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_262 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_427 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1539__B _1539_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1600__A2 _1256_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1274__B _1273_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_159 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_310 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1667__A2 _1608_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_259 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_207 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_74 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_387 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_421 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_62 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_402 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_262 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_95 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1052__B1 _1051_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_152 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1355__B2 SCAN_IN[18] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_137 VSS VDD sky130_fd_sc_hd__decap_6
X_1203_ _1202_/Y _1434_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_26_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_77_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_310 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1865__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_354 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_65_343 VSS VDD sky130_fd_sc_hd__decap_4
X_1134_ _1131_/X _1123_/X _1133_/Y _1728_/A VSS VDD sky130_fd_sc_hd__a21o_4
X_1065_ _1065_/A _1084_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_18_292 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_240 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1359__B SCAN_IN[19] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1043__B1 _1042_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1898_ _1898_/D _1092_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_68_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_18 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_339 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_107 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1822__B _1821_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1649__A2 _1646_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_192 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_302 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_398 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_207 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_357 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_224 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_240 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_262 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_257 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__B1 _1257_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_268 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_32 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_457 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_279 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1716__C _1716_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_435 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1888__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_140 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1451__C _1386_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_354 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_376 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_357 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_335 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1273__B1 _1094_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_295 VSS VDD sky130_fd_sc_hd__decap_6
X_1821_ _1716_/A _1821_/B _1821_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1257__A2_N _1256_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_276 VSS VDD sky130_fd_sc_hd__fill_2
X_1752_ _1753_/A _1745_/X _1752_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1195__A _1897_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1683_ _1653_/X _1674_/X _1682_/Y SCAN_IN[21] _1575_/Y _1683_/X VSS VDD sky130_fd_sc_hd__a32o_4
XANTENNA__1328__B2 _1327_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_398 VSS VDD sky130_fd_sc_hd__decap_8
X_1117_ _1114_/X _1104_/X _1117_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_65_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_357 VSS VDD sky130_fd_sc_hd__fill_1
X_1048_ _0976_/A _1037_/Y _1048_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_21_221 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1264__B1 _1261_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_243 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_0_125 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1833__A _1833_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_43 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_324 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_154 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_243 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_36 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1743__A _1743_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_107 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1462__B _1462_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1874__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_184 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_195 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1903__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_379 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_198 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1797__A1 _1719_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_390 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1549__A1 _1587_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1804_ _1803_/C _1804_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1549__B2 _1548_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1735_ _1737_/A _1751_/B _1735_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_7_291 VSS VDD sky130_fd_sc_hd__decap_3
X_1666_ _1347_/Y _1630_/A _1664_/Y _1665_/X _1676_/A VSS VDD sky130_fd_sc_hd__a211o_4
X_1597_ _1597_/A _1584_/X _1596_/Y _1597_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1075__D _1075_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1653__A SCAN_IN[20] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1721__A1 _1718_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_132 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1485__B1 _1478_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_195 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1788__B2 _1794_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1788__A1 _1719_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_23 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1828__A _1798_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_11 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_44 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_1_412 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_434 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1712__B2 _1711_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_140 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_324 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_184 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_121 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_96 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_357 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_143 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_44_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_316 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_71_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_51 VSS VDD sky130_fd_sc_hd__fill_2
X_1520_ _1359_/A _1520_/B _1523_/B VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1400__B1 _1399_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1451_ _1451_/A _1383_/B _1386_/C _1451_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_1382_ _1382_/A _1386_/C VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_67_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_327 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_102 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_clk_0_48_A clkbuf_0_clk_0_48/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1367__B _1345_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1718_ _1718_/A _1707_/Y _1718_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1649_ _1769_/A _1646_/B _1648_/Y _1649_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XANTENNA__1073__A2_N _1019_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1383__A _1218_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_460 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_110 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1830__B _1828_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_22 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_11 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_132 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_26_154 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_33 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_44 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_55 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_77 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_88 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_66 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_77 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_157 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_88 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_99 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0969__C1 _0968_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1558__A _1539_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_87 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1724__C _1716_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_26 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1697__B1 _1091_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_297 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_37 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_235 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_419 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1449__B1 _1196_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_110 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_17_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_293 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_433 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_319 VSS VDD sky130_fd_sc_hd__decap_12
X_0951_ _0951_/A _0945_/X _0951_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1621__B1 _1620_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1468__A _1525_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0975__A2 _0933_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_397 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_3 VSS VDD sky130_fd_sc_hd__decap_4
X_1503_ _1307_/A _1501_/X _1503_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1434_ _1434_/A _1379_/B _1434_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1365_ _1427_/A _1364_/Y _1347_/Y _1349_/B _1365_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1152__A2 _1143_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_419 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_249 VSS VDD sky130_fd_sc_hd__fill_2
X_1296_ _1228_/Y _1297_/B _1296_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_36_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_400 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_609 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_433 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1749__A1_N _1742_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_319 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1378__A _1378_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_190 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0966__A2 _1866_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_57 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1825__B _1822_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1391__A2 _1390_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_319 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1679__B1 _1663_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1841__A _1840_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_32 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1580__A2_N _1256_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_422 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1288__A _1285_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1603__B1 _1577_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_341 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_385 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_378 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1735__B _1751_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_69_319 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_50 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1751__A _1753_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1134__A2 _1123_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1150_ _1904_/Q _1143_/X _1150_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1470__B _1471_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1901__D _1901_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_441 VSS VDD sky130_fd_sc_hd__decap_8
X_1081_ _1081_/A _1078_/X _1081_/C _1080_/X _1081_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_37_249 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_400 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1198__A _1198_/A VSS VDD sky130_fd_sc_hd__diode_2
X_0934_ _1872_/Q _0933_/X _0934_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1373__A2 _1361_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1417_ _1261_/Y _1417_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_68_341 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1125__A2 _1118_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_396 VSS VDD sky130_fd_sc_hd__fill_1
X_1348_ _1239_/A _1349_/B VSS VDD sky130_fd_sc_hd__buf_1
X_1279_ _1279_/A _1264_/X _1278_/Y _1279_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_43_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_433 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_406 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1611__A1_N _1600_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_23 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_89 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1836__A _1833_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_330 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1329__B1_N _1328_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1571__A _1571_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_322 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_216 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_271 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_433 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_425 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1052__A1 _0991_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_182 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_69_116 VSS VDD sky130_fd_sc_hd__fill_2
X_1202_ _1146_/A _1202_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_19_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1133_ _1132_/X _1133_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1064_ _1923_/Q _1064_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_21_414 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_469 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1043__A1 _1040_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1897_ _1527_/X _1897_/Q _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_75_119 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_56_300 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_12 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_219 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_17_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_336 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1806__B1 _1788_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_225 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_414 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_258 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__B2 _1281_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1282__A1 _1202_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_269 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1566__A _1566_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_134 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_447 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_58_85 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_47_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_74_51 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_74_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_369 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1273__A1 _1096_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1273__B2 SCAN_IN[1] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_200 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_770 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_391 VSS VDD sky130_fd_sc_hd__decap_6
X_1820_ _1820_/A _1821_/B _1819_/Y _1820_/D _1820_/Y VSS VDD sky130_fd_sc_hd__nor4_4
XFILLER_30_266 VSS VDD sky130_fd_sc_hd__decap_8
X_1751_ _1753_/A _1751_/B _1751_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1476__A _1199_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1682_ _1675_/X _1681_/X _1673_/A _1682_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1916__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_333 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_314 VSS VDD sky130_fd_sc_hd__fill_2
X_1116_ _1115_/Y _1116_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1047_ _1041_/A _1046_/Y _1047_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1264__B2 _1262_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_233 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_277 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1386__A _1334_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1833__B _1831_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_137 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1302__A2_N _1264_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_355 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_163 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_314 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_188 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_215 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1296__A _1228_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1855__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1907__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_410 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_69_40 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_454 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1743__B _1694_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_73 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_62 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_67_406 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_141 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_133 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_325 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_62_177 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_328 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1797__A2 _1716_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1803_ _1803_/A _1797_/X _1803_/C _1803_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1549__A2 _1546_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1734_ _1734_/A _1716_/B _1716_/C _1734_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_1665_ _1364_/Y _1536_/A SCAN_IN[15] _1543_/B _1665_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
X_1596_ _1594_/Y _1596_/B _1596_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1653__B _1652_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1721__A2 _1719_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_417 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_66_450 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_163 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_100 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1485__A1 _1430_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1485__B2 _1484_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_38_185 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_369 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_339 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1878__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1788__A2 _1716_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1828__B _1824_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1880__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1844__A _1575_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_457 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_76_203 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1173__B1 _1107_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_258 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_236 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_39_98 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_55_42 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_328 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_199 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_380 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_8 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1400__A1 _1304_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1754__A _1754_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_7 VSS VDD sky130_fd_sc_hd__fill_2
X_1450_ _1405_/X _1442_/Y _1443_/X _1448_/X _1449_/X _1450_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XANTENNA__1904__D _1749_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1381_ _1376_/X _1383_/B VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1164__B1 _1119_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_420 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_339 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_188 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_114 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_50_169 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1367__C _1357_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1717_ _1719_/A _1695_/B _1717_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1664__A _1663_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1648_ _1602_/X _1647_/X _1602_/X _1647_/X _1648_/Y VSS VDD sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__1383__B _1383_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1579_ _1579_/A _1579_/B _1579_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1458__A1 _1421_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1830__C _1829_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_12 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_144 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_23 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_306 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_34 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_45 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_56 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_114 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_199 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_67 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_78 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1839__A _1833_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_89 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0969__B1 _0967_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_66 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1574__A _1571_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_210 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_232 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_1_265 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1697__A1 _1089_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1697__B2 _1566_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_64_239 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_57_280 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1449__A1 _1158_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_177 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_125 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_350 VSS VDD sky130_fd_sc_hd__decap_8
X_0950_ _0948_/A _0950_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1621__A1 SCAN_IN[0] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1468__B _1467_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1385__B1 _1379_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1502_ _1502_/A _1502_/B _1500_/Y _1501_/X _1502_/X VSS VDD sky130_fd_sc_hd__and4_4
X_1433_ _1405_/X _1427_/Y _1428_/X _1431_/Y _1432_/X _1880_/D VSS VDD sky130_fd_sc_hd__o32ai_4
XFILLER_49_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1364_ SCAN_IN[16] _1364_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1295_ _1257_/X _1281_/Y _1257_/X _1281_/Y _1297_/B VSS VDD sky130_fd_sc_hd__a2bb2oi_4
XFILLER_55_239 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_272 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_261 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_412 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1845__D1 _1820_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_445 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_423 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_158 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1659__A SCAN_IN[12] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_180 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1916__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_36 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1376__B1 _1375_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1394__A _1394_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1679__B2 _1665_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1679__A1 _1676_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_409 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_272 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_42_412 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_445 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_32 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_169 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1853__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_467 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1569__A _1575_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1603__A1 _1181_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1288__B _1287_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1603__B2 _1602_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_331 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_180 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_313 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_331 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_8 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_95 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_84 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1751__B _1751_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_397 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_375 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_453 VSS VDD sky130_fd_sc_hd__decap_4
X_1080_ _0964_/A _1866_/Q _0999_/X _0961_/B _1080_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_45_261 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_423 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_264 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1072__A2_N _1040_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_106 VSS VDD sky130_fd_sc_hd__fill_1
X_0933_ _1871_/Q _0932_/X _0933_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_9_184 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1373__A3 _1372_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1416_ _1349_/B _1408_/B _1408_/C _1416_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_68_353 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_92 VSS VDD sky130_fd_sc_hd__fill_2
X_1347_ SCAN_IN[15] _1347_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_28_206 VSS VDD sky130_fd_sc_hd__decap_8
X_1278_ _1276_/Y _1278_/B _1278_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1655__A2_N _1567_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_412 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_407 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_467 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_418 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_275 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_106 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_139 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1836__B _1834_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_139 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1571__B _1571_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_397 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_375 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_53 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_86 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_286 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1588__B1 _1587_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_150 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1052__A2 _1050_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0931__A _1869_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_194 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_143 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_12_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_176 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_7 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1762__A _1762_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_393 VSS VDD sky130_fd_sc_hd__decap_4
X_1201_ _1238_/B _1442_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_77_161 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_150 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1912__D _1823_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1132_ _1131_/X _1123_/X _1132_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_65_367 VSS VDD sky130_fd_sc_hd__decap_3
X_1063_ _0927_/X _1063_/B _1062_/X _1063_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_33_220 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_21_404 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_286 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_297 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1043__A2 _1041_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1896_ _1896_/D _1240_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_0_308 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_319 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_56_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_315 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1806__A1 _1795_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_79 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_215 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1282__A2 _1256_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1847__A _1847_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_78 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_415 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_404 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_3_168 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_426 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_459 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_59_172 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_97 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_59_194 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_315 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_304 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0926__A _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_389 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_197 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_337 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1273__A2 _1272_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_275 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_30_212 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_771 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _1790_/B _1716_/B _1716_/C _1750_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_30_289 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_7_441 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1476__B _1442_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1907__D _1907_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_452 VSS VDD sky130_fd_sc_hd__decap_12
X_1681_ _1674_/A _1679_/Y _1680_/Y _1654_/Y _1681_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1733__B1 _1728_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_345 VSS VDD sky130_fd_sc_hd__fill_1
X_1115_ _1114_/X _1115_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_38_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_53_337 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_0_71 VSS VDD sky130_fd_sc_hd__fill_1
X_1046_ _0976_/A _1044_/X _1045_/X _1046_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XFILLER_21_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_256 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_21_289 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1386__B _1383_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1879_ _1879_/D _1127_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA_clkbuf_1_1_0_clk_1_0_A clkbuf_0_clk_1_0/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__CTS_buf_1_32_A _CTS_buf_1_32/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_149 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1833__C _1832_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_23 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_323 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_29_345 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_29_367 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_71_123 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_71_112 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_56_175 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_337 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_348 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_71_167 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_71_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_52_370 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_44_99 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1577__A _1179_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_267 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_256 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_60_65 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_8_238 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1296__B _1297_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_52 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1743__C _1694_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_164 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_35_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_3 VSS VDD sky130_fd_sc_hd__decap_12
X_1802_ _1729_/A _1724_/A _1800_/Y _1801_/X _1803_/C VSS VDD sky130_fd_sc_hd__a211o_4
XPHY_590 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1733_ _1713_/X _1724_/Y _1726_/X _1728_/Y _1732_/X _1733_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
X_1664_ _1663_/X _1664_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1595_ _1587_/A SCAN_IN[2] _1585_/X _1585_/A SCAN_IN[3] _1596_/B VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_58_429 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_112 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_337 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1485__A2 _1427_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_145 VSS VDD sky130_fd_sc_hd__fill_1
X_1029_ _1028_/X _1029_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_14_36 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_14_69 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1397__A _1096_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1844__B _1844_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1173__A1 _1827_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_76_215 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_469 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1173__B2 _1172_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_462 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_57_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_315 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_54 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1100__A _1494_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_40_373 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_384 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1400__A2 _1397_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1164__A1 _1820_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1380_ _1897_/Q _1384_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1164__B2 _1163_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1770__A _1771_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_226 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_270 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1920__D _1848_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_123 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_50_137 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1367__D _1366_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1716_ _1716_/A _1716_/B _1716_/C _1716_/Y VSS VDD sky130_fd_sc_hd__nor3_4
X_1647_ _1772_/A SCAN_IN[9] _1577_/X _1647_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_6_81 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1900__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1383__C _1386_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_215 VSS VDD sky130_fd_sc_hd__fill_2
X_1578_ _1760_/A _1578_/B _1578_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1680__A _1655_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_218 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_410 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1458__A2 _1456_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1830__D _1827_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_454 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_13 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_318 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_35 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_46 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_24 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_57 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_68 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_79 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_351 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0969__A1 _0964_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1839__B _1837_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1441__A1_N _1434_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_56 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_78 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1574__B _1571_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_3 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_2_17 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_49_204 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1697__A2 _1696_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_215 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1449__A2 _1401_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_45_410 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_123 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_432 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_402 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0934__A _1872_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1621__A2 _1619_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_322 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1468__C _1468_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_388 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1385__A1 _1196_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1385__B2 _1384_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1915__D _1833_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1501_ _1216_/Y _1498_/X _1501_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1432_ _1140_/X _1412_/X _1196_/X _1432_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1868__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_1363_ _1894_/Q _1675_/A _1240_/B _1346_/Y _1366_/C VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_55_207 VSS VDD sky130_fd_sc_hd__decap_12
X_1294_ _1238_/B _1322_/B _1321_/A VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_36_410 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1005__A _1005_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_292 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1845__C1 _1844_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_295 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1659__B _1658_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1073__B1 _1868_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1675__A _1675_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1376__A1 SCAN_IN[21] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1394__B _1383_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1679__A2 _1669_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_421 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_432 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_251 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_104 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_52_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_457 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1569__B _1569_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_44 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_52_88 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1603__A2 _1577_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1893__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1585__A _1585_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_30 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0929__A _1865_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_229 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_276 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_20_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_170 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_192 VSS VDD sky130_fd_sc_hd__fill_2
X_0932_ _1870_/Q _0931_/X _0932_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1495__A _1492_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_3 VSS VDD sky130_fd_sc_hd__decap_8
X_1415_ _1405_/X _1408_/Y _1409_/X _1413_/Y _1414_/X _1415_/Y VSS VDD sky130_fd_sc_hd__o32ai_4
XFILLER_68_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_82 VSS VDD sky130_fd_sc_hd__decap_4
X_1346_ SCAN_IN[20] _1346_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_68_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_376 VSS VDD sky130_fd_sc_hd__fill_2
X_1277_ _1268_/A SCAN_IN[2] _1266_/X _1114_/X SCAN_IN[3] _1278_/B VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_24_402 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_408 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_243 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_419 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1836__C _1836_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_306 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_3_328 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_7 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_59_343 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_11 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_402 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_99 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1285__B1 _1249_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_42_254 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_276 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1588__A1 _1587_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1588__B2 SCAN_IN[2] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0931__B _0930_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_166 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1762__B _1762_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_140 VSS VDD sky130_fd_sc_hd__fill_2
X_1200_ _1165_/A _1200_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_77_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_335 VSS VDD sky130_fd_sc_hd__fill_2
X_1131_ _1583_/A _1131_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1906__CLK _1924_/Q VSS VDD sky130_fd_sc_hd__diode_2
X_1062_ _1061_/A _1061_/B _1062_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_18_251 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_254 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_449 VSS VDD sky130_fd_sc_hd__decap_12
X_1895_ _1895_/D _1240_/B _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_1_0_0_clk_1_0_A clkbuf_0_clk_1_0/X VSS VDD sky130_fd_sc_hd__diode_2
X_1329_ _1460_/A _1326_/B _1328_/Y _1329_/Y VSS VDD sky130_fd_sc_hd__a21boi_4
XFILLER_17_47 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1267__B1 _1266_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1806__A2 _1787_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_216 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_449 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_46 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1847__B _1847_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_184 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_176 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_75 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1103__A _1268_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_243 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_772 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0942__A _0942_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_11_460 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_7_464 VSS VDD sky130_fd_sc_hd__decap_6
X_1680_ _1655_/X _1680_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1733__B2 _1732_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1733__A1 _1713_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1923__D BB_IN VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_24_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_65_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_324 VSS VDD sky130_fd_sc_hd__fill_1
X_1114_ _1114_/A _1114_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_165 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_368 VSS VDD sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clk_0_48 clkbuf_0_clk_0_48/X _1924_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1925__RESET_B RESET_N VSS VDD sky130_fd_sc_hd__diode_2
X_1045_ _0976_/A _1044_/X _1045_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_0_94 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1013__A _0964_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_81 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_92 VSS VDD sky130_fd_sc_hd__decap_4
X_1878_ _1415_/Y _1114_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1386__C _1386_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_106 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1833__D _1827_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_302 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1488__B1 _1486_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_379 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_135 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_202 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_44_67 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_382 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_12_213 VSS VDD sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk_1_0 _CTS_root/X clkbuf_0_clk_1_0/X VSS VDD sky130_fd_sc_hd__clkbuf_16
XANTENNA__1577__B _1577_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_206 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1593__A _1593_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_31 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_79_246 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_67_419 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0937__A _1874_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_110 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_47_121 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1479__B1 _1245_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_176 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_62_146 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1768__A _1768_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1651__B1 _1777_/C VSS VDD sky130_fd_sc_hd__diode_2
X_1801_ _1737_/A _1734_/A _1131_/X _1543_/B _1801_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XPHY_580 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1918__D _1843_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1732_ _1727_/X _1731_/X _1529_/X _1732_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1403__B1 _1402_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_283 VSS VDD sky130_fd_sc_hd__fill_2
X_1663_ _1662_/X _1663_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1594_ _1594_/A _1589_/Y _1614_/A _1594_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_38_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_327 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_390 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_168 VSS VDD sky130_fd_sc_hd__decap_6
X_1028_ _0999_/X _0968_/A _1019_/Y _1028_/D _1028_/X VSS VDD sky130_fd_sc_hd__or4_4
XANTENNA__1642__B1 _1743_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_15 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_48 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1397__B _1098_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_30_25 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_30_36 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_426 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1173__A2 _1168_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_408 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_419 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_110 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_411 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1330__C1 _1329_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_165 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_55_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_135 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1633__B1 _1596_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_76 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_396 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_67_205 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1164__A2 _1158_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1770__B _1751_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_238 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1639__A1_N _1580_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_293 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_444 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_319 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1498__A _1217_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1624__B1 _1614_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_149 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_385 VSS VDD sky130_fd_sc_hd__fill_2
X_1715_ _1690_/A _1716_/C VSS VDD sky130_fd_sc_hd__buf_1
X_1646_ _1769_/A _1646_/B _1646_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_6_93 VSS VDD sky130_fd_sc_hd__decap_8
X_1577_ _1179_/Y _1577_/B _1577_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_58_238 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_260 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_26_102 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_444 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_433 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_14 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_36 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_47 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_58 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_69 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_127 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1615__B1 _1614_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1201__A _1238_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1839__C _1839_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_385 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0969__A2 _0959_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_245 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_1_278 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_49_238 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_32 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_49_249 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_208 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_455 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_263 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_414 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0934__B _0933_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1606__B1 _1578_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_396 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0950__A _0948_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1385__A2 _1244_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1500_ _1216_/Y _1498_/X _1500_/Y VSS VDD sky130_fd_sc_hd__nand2_4
X_1431_ _1429_/X _1430_/X _1412_/X _1431_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1781__A _1720_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1362_ SCAN_IN[19] _1675_/A VSS VDD sky130_fd_sc_hd__inv_8
X_1293_ _1282_/X _1292_/X _1282_/X _1292_/X _1322_/B VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_219 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1845__B1 _1502_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_127 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1021__A _1019_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1073__B2 _1019_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_160 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1675__B _1759_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1376__A2 _1525_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1394__C _1386_/C VSS VDD sky130_fd_sc_hd__diode_2
X_1629_ _1596_/Y _1584_/X _1596_/Y _1584_/X _1629_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1691__A _1547_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1679__A3 _1678_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_46_219 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_296 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_116 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_14_138 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1569__C _1569_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_344 VSS VDD sky130_fd_sc_hd__fill_2
X_CTS_buf_1_32 _CTS_buf_1_32/A _CTS_buf_1_32/X VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1585__B SCAN_IN[3] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_326 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_337 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1862__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0929__B _1866_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_75 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_255 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_447 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_458 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_288 VSS VDD sky130_fd_sc_hd__decap_12
X_0931_ _1869_/Q _0930_/X _0931_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1776__A _1683_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_164 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_54_3 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_381 VSS VDD sky130_fd_sc_hd__fill_2
X_1414_ _1118_/X _1412_/X _1196_/X _1414_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_1345_ _1394_/A _1339_/Y _1342_/X _1344_/Y _1345_/X VSS VDD sky130_fd_sc_hd__a211o_4
XANTENNA__1016__A _0999_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1276_ _1276_/A _1270_/X _1276_/C _1276_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_36_252 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_51_233 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_409 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1046__A1 _0976_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1686__A _1686_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_48 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1836__D _1827_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_318 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_59_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_355 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_47_78 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1809__B1 _1792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_230 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1285__B2 _1284_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1285__A1 _1176_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_263 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_296 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_42_266 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1596__A _1594_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1588__A2 _1269_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1858__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_101 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_123 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_69_108 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1762__C _1762_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_303 VSS VDD sky130_fd_sc_hd__fill_2
X_1130_ _1127_/X _1117_/X _1129_/Y _1130_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_77_196 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_347 VSS VDD sky130_fd_sc_hd__fill_1
X_1061_ _1061_/A _1061_/B _1063_/B VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_18_263 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_296 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_428 VSS VDD sky130_fd_sc_hd__decap_4
X_1894_ _1521_/X _1894_/Q _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_68_141 VSS VDD sky130_fd_sc_hd__decap_12
X_1328_ _1284_/X _1327_/X _1284_/X _1327_/X _1328_/Y VSS VDD sky130_fd_sc_hd__a2bb2oi_4
XFILLER_71_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_17_26 VSS VDD sky130_fd_sc_hd__decap_6
X_1259_ _1259_/A SCAN_IN[5] _1259_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_71_339 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_328 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1267__A1 _1115_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_59 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_206 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_239 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_266 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_33_14 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_152 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_141 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_58_77 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_58_66 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_122 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_144 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_43 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_32 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_98 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_350 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_762 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1733__A2 _1724_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1194__B1 _1193_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_450 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_3 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_53_306 VSS VDD sky130_fd_sc_hd__decap_6
X_1113_ _1100_/X _1113_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_65_188 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_65_177 VSS VDD sky130_fd_sc_hd__fill_2
X_1044_ _1040_/X _1034_/X _1044_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1013__B _1013_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_71 VSS VDD sky130_fd_sc_hd__decap_8
X_1877_ _1404_/X _1268_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_69_461 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1488__B2 _1487_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1488__A1 _1452_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_133 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1204__A _1238_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_328 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_44_24 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_52_394 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_60_56 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_20_280 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_5_18 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_402 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0937__B _0935_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1479__B2 _1218_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1479__A1 _1097_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1114__A _1114_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_306 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_188 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_47_199 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_62_158 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1224__A1_N _1115_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1768__B _1767_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_70_180 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1651__A1 _1777_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_383 VSS VDD sky130_fd_sc_hd__decap_4
X_1800_ _1800_/A _1800_/Y VSS VDD sky130_fd_sc_hd__inv_8
XPHY_570 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ _1729_/A _1719_/X _1730_/Y _1731_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1403__A1 _1106_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_262 VSS VDD sky130_fd_sc_hd__decap_4
X_1662_ SCAN_IN[16] _1798_/B _1662_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1593_ _1593_/A _1614_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1024__A _1023_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1027_ _1023_/Y _1068_/B _1028_/D VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1642__A1 _1790_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1642__B2 _1639_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1397__C _1397_/C VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1919__CLK _1920_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1694__A _1694_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_416 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1158__B1 _1157_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_68 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_55_34 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1330__B1 _1326_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_456 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1887__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_361 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1633__A1 _1729_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_0_32_A _CTS_buf_1_32/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_55 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_71_33 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1633__B2 _1584_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_99 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1109__A _1108_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_243 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1149__B1 _1148_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0948__A _0948_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_67_217 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_261 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_35_136 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1779__A _1778_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1624__A1 _1593_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_372 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1498__B _1219_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_331 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_364 VSS VDD sky130_fd_sc_hd__fill_2
X_1714_ _1689_/A _1716_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_6_50 VSS VDD sky130_fd_sc_hd__decap_8
X_1645_ _1608_/X _1612_/X _1643_/Y _1759_/A _1608_/B _1646_/B VSS VDD sky130_fd_sc_hd__a32o_4
XANTENNA__1019__A _0963_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1576_ _1575_/Y _1777_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_58_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1560__B1 _1559_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1312__B1 _1274_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1689__A _1689_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_467 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_309 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_37 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_48 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_59 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_59 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_41_106 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1615__A1 _1587_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_320 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_180 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_191 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1839__D _1827_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1891__CLK _1887_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_257 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1551__B1 _1549_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_22 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_77 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_66_66 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_55 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_17_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_423 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1599__A _1597_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_17_169 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_45_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_106 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1606__A1 _1169_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_70 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1385__A3 _1245_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1430_ _1430_/A _1422_/X _1430_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1781__B _1781_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1361_ _1361_/A SCAN_IN[16] _1361_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_0_290 VSS VDD sky130_fd_sc_hd__decap_12
X_1292_ _1157_/A SCAN_IN[7] _1254_/X _1292_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_36_434 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_36_445 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1845__A1 _1777_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_253 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_404 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_51_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_139 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1021__B _1018_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_172 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_194 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_17 VSS VDD sky130_fd_sc_hd__fill_2
X_1628_ _1544_/A _1716_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1691__B _1694_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1559_ _1905_/Q _1557_/Y _1539_/X _1169_/X _1558_/X _1559_/Y VSS VDD sky130_fd_sc_hd__a32oi_4
XFILLER_42_404 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_54_286 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_264 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1212__A _1211_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1569__D _1568_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_323 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_312 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_194 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0929__C _1867_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_45_231 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_242 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1122__A _1585_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_404 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_275 VSS VDD sky130_fd_sc_hd__fill_2
X_0930_ _1868_/Q _0929_/X _0930_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__0961__A _0959_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_121 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_9_176 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_42_90 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1792__A _1792_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1413_ _1410_/X _1411_/X _1412_/X _1413_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1919__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_323 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_3_62 VSS VDD sky130_fd_sc_hd__decap_3
X_1344_ _1343_/X _1344_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1275_ _1094_/X SCAN_IN[1] _1274_/X _1276_/C VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1016__B _1015_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_212 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1032__A _0998_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_437 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1046__A2 _1044_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_38 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__CTS_buf_1_48_A _CTS_buf_1_0/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1207__A _1352_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1852__D _1852_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_334 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_378 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_367 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_24 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_337 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_326 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1809__A1 _1803_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1809__B2 _1790_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1285__A2 _1577_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_275 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_67 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_34 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1562__A1_N _1812_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_223 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_78 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_429 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1596__B _1596_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_135 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_71 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_6_146 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_352 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1117__A _1114_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0956__A _0955_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_315 VSS VDD sky130_fd_sc_hd__decap_12
X_1060_ _1058_/A _1060_/B _1037_/Y _1061_/B VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_33_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_278 VSS VDD sky130_fd_sc_hd__fill_2
X_1893_ _1893_/D _1238_/B _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1027__A _1023_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_186 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_56_337 VSS VDD sky130_fd_sc_hd__decap_12
X_1327_ _1463_/A SCAN_IN[9] _1249_/X _1327_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_1258_ SCAN_IN[5] _1258_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_17_16 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1267__A2 _1265_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1189_ _1885_/Q _1189_/Y VSS VDD sky130_fd_sc_hd__inv_8
XPHY_207 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_418 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_229 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_105 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_116 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_138 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_58_12 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_315 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_189 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_245 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_278 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_763 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_774 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_422 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_400 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1194__A1 _1113_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1733__A3 _1726_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1902__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_123 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_65_112 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_337 VSS VDD sky130_fd_sc_hd__fill_2
X_1112_ _1064_/X _1106_/X _1107_/X _1111_/X _1112_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_53_318 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_30 VSS VDD sky130_fd_sc_hd__fill_1
X_1043_ _1040_/X _1041_/X _1042_/Y _1043_/X VSS VDD sky130_fd_sc_hd__o21a_4
XFILLER_0_74 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_63 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1310__A _1273_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_237 VSS VDD sky130_fd_sc_hd__decap_6
X_1876_ _1392_/X _1094_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1488__A2 _1451_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_315 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_29_326 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_337 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_145 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_359 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_115 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_104 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_44_318 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_36 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_12_248 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_270 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_69_11 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_66 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_69_44 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_79_226 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_69_88 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1479__A2 _1217_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_454 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_47_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_47_145 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_340 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1651__A2 _1605_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_571 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_91 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_593 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ _1730_/A _1730_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_11_281 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_11_270 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1403__A2 _1388_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1661_ _1346_/Y _1569_/B _1657_/X _1659_/X _1660_/X _1661_/X VSS VDD sky130_fd_sc_hd__a2111o_4
X_1592_ _1091_/A SCAN_IN[1] _1591_/X _1593_/A VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_78_281 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_410 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_78_292 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_53_104 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1024__B _1022_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_26_318 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_38_167 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_148 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_189 VSS VDD sky130_fd_sc_hd__decap_4
X_1026_ _1014_/A _1024_/Y _1025_/X _1855_/D VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1642__A2 _1611_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1040__A _0980_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1694__B _1694_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1859_ _1859_/D _0973_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1158__A1 _1443_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_428 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1860__D _1860_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_69_292 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_123 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1215__A _1215_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1330__A1 _1247_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_178 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_351 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_384 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1633__A2 _1263_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1856__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_71_67 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_398 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_211 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1109__B _1090_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1149__A1 _1147_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_60 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_93 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0948__B _0947_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_443 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0964__A _0964_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1779__B _1772_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_170 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1624__A2 _1589_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_343 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1795__A _1089_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_376 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_77_3 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_390 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _1703_/A _1713_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_6_84 VSS VDD sky130_fd_sc_hd__fill_2
X_1644_ _1608_/A _1759_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1575_ _1575_/A _1575_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1560__A1 _1533_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1035__A _1011_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_421 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1312__A1 _1219_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1270__A1_N _1304_/A VSS VDD sky130_fd_sc_hd__diode_2
XPHY_16 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_38 VSS VDD sky130_fd_sc_hd__decap_3
X_1009_ _1000_/Y _1008_/X _0991_/Y _0995_/A _1009_/X VSS VDD sky130_fd_sc_hd__a211o_4
XPHY_49 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_170 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_41_118 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1615__A2 _1269_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_332 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_398 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_41_48 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_59 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1855__D _1855_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_225 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_236 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1551__B2 _1550_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1551__A1 _1718_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_89 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_57_284 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_72_243 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1599__B _1598_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_276 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_332 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_181 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1606__A2 SCAN_IN[8] VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_376 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_15_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1869__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_358 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_336 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_81 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0959__A _1865_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1781__C _1780_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1360_ _1359_/X _1366_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_0_280 VSS VDD sky130_fd_sc_hd__decap_4
X_1291_ _1283_/X _1290_/Y _1291_/X VSS VDD sky130_fd_sc_hd__xor2_4
XANTENNA__1909__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_251 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_63_221 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_210 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_424 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1845__A2 _1842_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_457 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_276 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_416 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_184 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1230__B1 _1166_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1627_ _1805_/B _1617_/Y _1625_/Y _1626_/Y _1627_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1691__C _1694_/C VSS VDD sky130_fd_sc_hd__diode_2
X_1558_ _1539_/B _1558_/X VSS VDD sky130_fd_sc_hd__buf_1
X_1489_ _1166_/A _1359_/A _1176_/A _1460_/A _1489_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_15 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_54_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_427 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_335 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_6_317 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_55 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_357 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_402 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_457 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_265 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_60_268 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0961__B _0961_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_13_184 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_42_80 VSS VDD sky130_fd_sc_hd__decap_8
X_1412_ _1237_/A _1412_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_3_52 VSS VDD sky130_fd_sc_hd__decap_4
X_1343_ _1342_/A _1341_/Y _1394_/A _1339_/Y _1343_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_68_357 VSS VDD sky130_fd_sc_hd__fill_1
X_1274_ _1274_/A _1273_/X _1274_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1016__C _1011_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1881__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_36_210 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_416 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_265 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_36_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_279 VSS VDD sky130_fd_sc_hd__fill_1
X_0989_ _0992_/A _0991_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_74_349 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1809__A2 _1808_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1223__A _1216_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_202 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_57 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_408 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_10_154 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_50 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_158 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_83 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0953__C1 _0952_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1117__B _1104_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_165 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_65_327 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1133__A _1132_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_232 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_371 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_276 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_33_202 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_393 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0972__A _0971_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1681__B1 _1680_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_21_419 VSS VDD sky130_fd_sc_hd__decap_4
X_1892_ _1515_/X _1198_/A _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1433__B1 _1431_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1308__A _1211_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1027__B _1068_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_154 VSS VDD sky130_fd_sc_hd__decap_12
X_1326_ _1460_/A _1326_/B _1326_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XFILLER_56_316 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1325__B1_N _1324_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_56_349 VSS VDD sky130_fd_sc_hd__decap_12
X_1257_ _1202_/Y _1256_/X _1202_/Y _1255_/Y _1257_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_319 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_64_371 VSS VDD sky130_fd_sc_hd__fill_2
X_1188_ _1771_/A _1171_/Y _1908_/Q _1778_/A _1182_/X _1188_/X VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_24_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1672__B1 SCAN_IN[13] VSS VDD sky130_fd_sc_hd__diode_2
XPHY_219 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_38 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_441 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1424__B1 _1423_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1218__A _1218_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1863__D _1113_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_102 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_59_176 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_198 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_74_168 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_62_319 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_308 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_55_382 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_224 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_235 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_720 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 VSS VDD sky130_fd_sc_hd__decap_12
XPHY_753 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_441 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1415__B1 _1413_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_71 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1128__A _1127_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1194__A2 _1188_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_7 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__0967__A _0968_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_194 VSS VDD sky130_fd_sc_hd__decap_12
X_1111_ _1108_/X _1090_/X _1110_/Y _1111_/X VSS VDD sky130_fd_sc_hd__a21o_4
XFILLER_65_157 VSS VDD sky130_fd_sc_hd__fill_2
X_1042_ _1040_/X _1041_/X _1032_/X _1042_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XANTENNA__1798__A _1736_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_385 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_205 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_290 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_21_249 VSS VDD sky130_fd_sc_hd__fill_1
X_1875_ _1875_/D _1271_/A _1847_/X _1923_/Q VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1038__A _0950_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_102 VSS VDD sky130_fd_sc_hd__decap_12
X_1309_ _1276_/C _1270_/X _1276_/C _1270_/X _1309_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_371 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1645__B1 _1759_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1501__A _1216_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_205 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1858__D _1043_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_69 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_23 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_249 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_79_238 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_79_216 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_75_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_400 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_47_102 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_75_466 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_371 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1636__B1 _1724_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1411__A _1116_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_561 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_81 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_550 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_242 VSS VDD sky130_fd_sc_hd__fill_2
X_1660_ SCAN_IN[13] _1794_/B _1660_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1591_ _1092_/A SCAN_IN[0] _1590_/X _1591_/X VSS VDD sky130_fd_sc_hd__and3_4
XFILLER_7_297 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_38_179 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_53_116 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1627__B1 _1625_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1321__A _1321_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1025_ _1023_/Y _1022_/B _1025_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_34_330 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_341 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1328__A2_N _1327_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1694__C _1694_/C VSS VDD sky130_fd_sc_hd__diode_2
X_1858_ _1043_/X _0978_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1789_ _1789_/A _1786_/Y _1787_/X _1788_/X _1789_/X VSS VDD sky130_fd_sc_hd__and4_4
XFILLER_1_407 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1158__A2 _1148_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_411 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_400 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_444 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_135 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1330__A2 _1288_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_58 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_127 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_171 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_25_396 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_333 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_40_355 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_377 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_388 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1896__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_clk_0_48 clkbuf_0_clk_0_48/X _1923_/CLK VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1149__A2 _1139_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_451 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1406__A _1376_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_81 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_455 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_75_274 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_436 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1141__A _1903_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_341 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_385 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_91 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0980__A _0980_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_322 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_43_182 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_193 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1795__B _1658_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_380 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1712_ _1701_/X _1703_/X _1709_/X _1711_/X _1712_/X VSS VDD sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1793__C1 _1792_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1643_ _1637_/X _1641_/Y _1642_/Y _1643_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_6_63 VSS VDD sky130_fd_sc_hd__decap_12
X_1574_ _1571_/A _1571_/B _1574_/X VSS VDD sky130_fd_sc_hd__and2_4
XANTENNA__1316__A _1309_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1560__A2 _1537_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_400 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1848__B1 _1064_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1312__A2 _1311_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_285 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_66_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_425 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_17 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_28 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_190 VSS VDD sky130_fd_sc_hd__fill_2
X_1008_ _1001_/Y _1006_/X _0977_/D _1007_/Y _1008_/X VSS VDD sky130_fd_sc_hd__a211o_4
XPHY_39 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_28 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_22_311 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_22_366 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1871__D _1871_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1551__A2 _1794_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1205__A2_N _1442_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_49_219 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_296 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_45_436 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_299 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_60_439 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_311 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_388 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_56_9 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1136__A _1100_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1290_ _1165_/A SCAN_IN[8] _1252_/X _1290_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
XFILLER_48_263 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_56_90 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_16_171 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_193 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_31_141 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1230__B2 _1516_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1230__A1 _1157_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_392 VSS VDD sky130_fd_sc_hd__decap_4
X_1626_ _1623_/X _1624_/Y _1626_/Y VSS VDD sky130_fd_sc_hd__nor2_4
X_1557_ _1638_/A _1557_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1488_ _1452_/A _1451_/A _1486_/Y _1487_/X _1488_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_27_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_27 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_39_285 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_54_244 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_27_436 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_39_296 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_15 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1866__D _1112_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_10_358 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_307 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_329 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_34 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_211 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_60 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_428 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_26_82 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_93 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1712__A2_N _1703_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_123 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_13_174 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_156 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_145 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_196 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_373 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_5_362 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0971__B1 _0963_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1411_ _1116_/X _1398_/X _1411_/X VSS VDD sky130_fd_sc_hd__or2_4
X_1342_ _1342_/A _1341_/Y _1342_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1273_ _1096_/Y _1272_/Y _1094_/X SCAN_IN[1] _1273_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1299__A1_N _1279_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_24_428 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_36_299 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_450 VSS VDD sky130_fd_sc_hd__decap_8
X_0988_ _1860_/Q _0992_/A VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__0962__B1 _0929_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_303 VSS VDD sky130_fd_sc_hd__fill_2
X_1609_ _1609_/A _1790_/B VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_59_347 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1504__A _1307_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_59 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_27_211 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_222 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_417 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_428 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_299 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_0_0_A _CTS_buf_1_0/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_104 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_332 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__0953__B1 _1005_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_2_387 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_398 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_77_144 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_77_188 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_177 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_339 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_65_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_211 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1130__B1 _1129_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_383 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_288 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_214 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_236 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1681__B2 _1654_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1681__A1 _1674_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_14_450 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_269 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_80 VSS VDD sky130_fd_sc_hd__fill_2
X_1891_ _1512_/X _1238_/D _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1433__A1 _1405_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1433__B2 _1432_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1308__B _1302_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_122 VSS VDD sky130_fd_sc_hd__fill_1
X_1325_ _1451_/A _1291_/X _1324_/X _1326_/B VSS VDD sky130_fd_sc_hd__a21bo_4
XFILLER_68_166 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1324__A _1321_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1256_ _1255_/Y _1256_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_64_361 VSS VDD sky130_fd_sc_hd__decap_8
X_1187_ _1812_/A _1778_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_24_225 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1672__B2 _1794_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1672__A1 _1341_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_209 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_269 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_28 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_20_431 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1424__A1 _1417_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_32_280 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_453 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1188__B1 _1778_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_58_36 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_114 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_47_306 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_136 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_47_339 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1112__B1 _1107_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_79 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_70_320 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_0_48_A _CTS_buf_1_48/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_710 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_269 VSS VDD sky130_fd_sc_hd__decap_6
XPHY_754 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1415__A1 _1405_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1415__B2 _1414_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_413 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_23_50 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_94 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1871__CLK _1886_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1409__A _1116_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1128__B _1117_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0967__B _0968_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1110_ _1110_/A _1110_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_38_328 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_65_136 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_10 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_80 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_65_169 VSS VDD sky130_fd_sc_hd__fill_2
X_1041_ _1041_/A _1034_/X _1041_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_0_32 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0983__A _0983_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_350 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_73_180 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1798__B _1798_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_342 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_331 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_217 VSS VDD sky130_fd_sc_hd__decap_4
X_1874_ _1194_/Y _1874_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1319__A _1319_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1038__B _1037_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1590__B1 _1091_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1054__A _0991_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_114 VSS VDD sky130_fd_sc_hd__decap_3
X_1308_ _1211_/Y _1302_/Y _1308_/X VSS VDD sky130_fd_sc_hd__and2_4
X_1239_ _1239_/A _1214_/A _1216_/A _1217_/A _1239_/X VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_71_139 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1645__A1 _1608_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_361 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_44_16 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1645__B2 _1608_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_342 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1501__B _1498_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_60_15 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1894__CLK _1911_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1874__D _1194_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1229__A _1228_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_79 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_434 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_50 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_62_139 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1636__A1 _1734_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_72 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_361 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_383 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1636__B2 _1629_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_191 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1411__B _1398_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_43_364 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_562 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_232 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_254 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1139__A _1138_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1590_ _1091_/Y _1272_/Y _1091_/A SCAN_IN[1] _1590_/X VSS VDD sky130_fd_sc_hd__o22a_4
XFILLER_7_287 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0978__A _0978_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_250 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_66_434 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_3 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_66_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_38_158 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_53_128 VSS VDD sky130_fd_sc_hd__fill_2
X_1024_ _1023_/Y _1022_/B _1024_/Y VSS VDD sky130_fd_sc_hd__nand2_4
XANTENNA__1627__A1 _1805_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1627__B2 _1626_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1321__B _1296_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_191 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1049__A _1032_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1857_ _1857_/D _0946_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_30_29 VSS VDD sky130_fd_sc_hd__fill_2
X_1788_ _1719_/A _1716_/A _1108_/X _1794_/B _1788_/X VSS VDD sky130_fd_sc_hd__o22a_4
XANTENNA__1482__A2_N _1216_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1563__B1 _1181_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1315__B1 _1216_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__CTS_buf_1_16_A _CTS_buf_1_32/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_26 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1512__A _1506_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_72_448 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1869__D _1145_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_320 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_37_180 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_44_139 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_364 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_71_47 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_183 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_40_312 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_40_323 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_202 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_4_235 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1554__B1 _1551_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_84 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_430 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1306__B1 _1276_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_463 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_412 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_253 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_75_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_48_467 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_75_297 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_63_426 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1422__A _1417_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_106 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_16_320 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_43_150 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0980__B _0979_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_370 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_381 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1711_ _1111_/X _1696_/X _1762_/A _1711_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1793__B1 _1790_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1642_ _1790_/B _1611_/X _1743_/A _1639_/X _1642_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
XFILLER_6_42 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_6_75 VSS VDD sky130_fd_sc_hd__decap_6
X_1573_ _1698_/A _1573_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1316__B _1314_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1560__A3 _1540_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1848__A1 _1713_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_242 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_39_445 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_456 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_106 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_128 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1332__A _1332_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_459 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_18 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_29 VSS VDD sky130_fd_sc_hd__decap_3
X_1007_ _0980_/A _0979_/X _1007_/C _1007_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XFILLER_22_389 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_41_28 VSS VDD sky130_fd_sc_hd__decap_6
X_1909_ _1909_/D _1547_/A _1847_/X _1911_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1784__B1 _1771_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1507__A _1212_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_36 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_66_58 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_57_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_212 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_201 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_404 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1242__A _1245_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_72_223 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_301 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_367 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_62 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_40_175 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1775__B1 _1773_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1527__B1 _1113_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1417__A _1261_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_459 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0991__A _0991_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_120 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_153 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1908__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1766__B1 _1688_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_382 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1230__A2 _1513_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1625_ _1623_/X _1624_/Y _1702_/A _1625_/Y VSS VDD sky130_fd_sc_hd__a21oi_4
X_1556_ _1904_/Q _1798_/B _1543_/X _1555_/X _1556_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
X_1487_ _1434_/A _1198_/X _1476_/X _1443_/A _1442_/A _1487_/X VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_39_220 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_242 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_253 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1062__A _1061_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_404 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_50_440 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_50_451 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_348 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_337 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1757__B1 _1529_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1882__D _1450_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1237__A _1237_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_415 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_437 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_459 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_45_245 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_204 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_60_226 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_60_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_259 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_9_113 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_41_462 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1748__B1 _1762_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_9_168 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_42_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1881__SET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_54_7 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_5_385 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1147__A _1147_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0947__B1_N _0932_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0971__B2 _0962_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0971__A1 _0955_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1410_ _1114_/X _1399_/Y _1410_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_68_337 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0986__A _0953_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_43 VSS VDD sky130_fd_sc_hd__fill_2
X_1341_ SCAN_IN[14] _1341_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1272_ SCAN_IN[1] _1272_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_36_256 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_51_237 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_51_259 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1739__B1 _1529_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0987_ _0983_/A _1061_/A VSS VDD sky130_fd_sc_hd__buf_1
X_1608_ _1608_/A _1608_/B _1608_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1057__A _1041_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0962__A1 _0958_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_315 VSS VDD sky130_fd_sc_hd__decap_12
X_1539_ _1169_/X _1539_/B _1539_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_74_318 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1504__B _1501_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_49 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_245 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_267 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1520__A _1359_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_27_278 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_42_215 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_42_226 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1877__D _1404_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_30 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_2_322 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0953__A1 _1068_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_77_123 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1130__A1 _1127_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_37_82 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1666__C1 _1665_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1430__A _1430_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1681__A2 _1679_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1433__A2 _1427_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1890_ _1890_/D _1239_/A _1847_/X _1887_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_45_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_68_112 VSS VDD sky130_fd_sc_hd__fill_2
X_1324_ _1321_/Y _1323_/Y _1324_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1605__A _1603_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1324__B _1323_/Y VSS VDD sky130_fd_sc_hd__diode_2
X_1255_ SCAN_IN[6] _1255_/Y VSS VDD sky130_fd_sc_hd__inv_8
X_1186_ _1186_/A _1812_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_24_215 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1340__A _1214_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1672__A2 _1544_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_18 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1424__A2 _1411_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1188__B2 _1182_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1188__A1 _1771_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_101 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_59_145 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_59_123 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_58_48 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1515__A _1506_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_156 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_74_148 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_74_47 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1112__A1 _1064_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1112__B2 _1111_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_711 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_332 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1250__A _1200_/Y VSS VDD sky130_fd_sc_hd__diode_2
XPHY_744 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_421 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1415__A2 _1408_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_23_40 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_62 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_7_436 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1409__B _1379_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_65_104 VSS VDD sky130_fd_sc_hd__fill_2
X_1040_ _0980_/A _1040_/X VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_0_44 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__0983__B _0937_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_362 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1160__A _1579_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_395 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_53 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_229 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1811__C1 _1810_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1873_ _1184_/Y _1873_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1319__B _1303_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1590__B2 SCAN_IN[1] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1590__A1 _1091_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1335__A SCAN_IN[12] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1054__B _1045_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_28_29 VSS VDD sky130_fd_sc_hd__fill_2
X_1307_ _1307_/A _1306_/Y _1307_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_56_159 VSS VDD sky130_fd_sc_hd__fill_2
X_1238_ _1894_/Q _1238_/B _1198_/A _1238_/D _1240_/C VSS VDD sky130_fd_sc_hd__or4_4
XFILLER_64_170 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_64_181 VSS VDD sky130_fd_sc_hd__fill_1
X_1169_ _1906_/Q _1169_/X VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1645__A2 _1612_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_332 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1070__A _1870_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1912__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_398 VSS VDD sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_clk_1_0 clkbuf_0_clk_1_0/X _CTS_buf_1_0/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XANTENNA__1802__C1 _1801_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_251 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1030__B1 _0998_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_218 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_69_69 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1890__D _1890_/D VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1245__A _1245_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1665__A2_N _1536_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_115 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_47_137 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_18_62 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_62_107 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_18_84 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1636__A2 _1634_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_181 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_395 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_70_140 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_70_184 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_552 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_387 VSS VDD sky130_fd_sc_hd__fill_1
XPHY_530 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_240 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_295 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_266 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1139__B _1128_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_50_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1155__A _1155_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_402 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_66_413 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_373 VSS VDD sky130_fd_sc_hd__decap_12
X_1023_ _0955_/A _1023_/Y VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_34_310 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1088__B1 _1085_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1627__A2 _1617_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_181 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_61_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_140 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1321__C _1320_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_61_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_34_398 VSS VDD sky130_fd_sc_hd__fill_2
X_1925_ BB_IN DATA_OUT RESET_N CLK_OUT VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1856_ _1031_/Y _0943_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1260__B1 _1259_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1787_ _1089_/X _1658_/X _1619_/X _1787_/X VSS VDD sky130_fd_sc_hd__o21a_4
XANTENNA__1049__B _1047_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1563__B2 _1608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1563__A1 _1186_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1065__A _1065_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_28 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1315__A1 _1309_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_284 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_438 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_55_38 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1079__B1 _0928_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1512__B _1502_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1861__CLK _1853_/CLK VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_52_151 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_376 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1885__D _1474_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_247 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1003__B1 _0971_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1554__B2 _1553_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1554__A1 _1131_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_221 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1306__B2 _1305_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_29_50 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1703__A _1703_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_63_416 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1422__B _1411_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_35_118 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_129 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_28_170 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_28_192 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1490__B1 _1488_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_398 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_31_335 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_162 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_184 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_360 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_1710_ _1688_/A _1762_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1793__A1 _1745_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1641_ _1743_/A _1639_/X _1640_/X _1641_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XFILLER_6_32 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__0989__A _0992_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1572_ _1571_/X _1698_/A VSS VDD sky130_fd_sc_hd__buf_1
XANTENNA__1560__A4 _1556_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1884__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_413 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1848__A2 _1813_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1613__A _1613_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_39_468 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_276 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_19 VSS VDD sky130_fd_sc_hd__decap_3
X_1006_ _0957_/A _1003_/Y _1004_/Y _1005_/Y _0952_/Y _1006_/X VSS VDD sky130_fd_sc_hd__a32o_4
XFILLER_34_140 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_162 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1481__B1 _1479_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_22_346 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_195 VSS VDD sky130_fd_sc_hd__decap_12
X_1908_ _1783_/Y _1908_/Q _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1233__B1 _1176_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1784__A1 _1763_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1784__B2 _1769_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1839_ _1833_/A _1837_/X _1839_/C _1827_/D _1839_/X VSS VDD sky130_fd_sc_hd__and4_4
XFILLER_1_206 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1507__B _1503_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_26 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_57_232 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1523__A _1333_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1242__B _1245_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_30 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_173 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_25_184 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_9_306 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_132 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_85 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_40_154 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1224__B1 _1127_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1775__A1 _1762_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1775__B2 _1774_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_62 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_31_95 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1527__A1 _1405_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_261 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_416 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_276 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_213 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_70 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_36_438 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_36_449 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_48_298 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_63_279 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0991__B _0990_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_16_140 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_72_80 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_3 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_190 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1766__A1 _1172_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_8_361 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1608__A _1608_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1230__A3 _1208_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1624_ _1593_/A _1589_/A _1614_/X _1624_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
X_1555_ _1736_/A _1543_/B _1554_/X _1555_/X VSS VDD sky130_fd_sc_hd__a21o_4
X_1486_ _1147_/A _1513_/A _1475_/X _1477_/Y _1485_/Y _1486_/Y VSS VDD sky130_fd_sc_hd__a2111oi_4
XFILLER_27_416 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_39_265 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_54_213 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1062__B _1061_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_42_408 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_132 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_316 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_10_305 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_22_154 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_10_327 VSS VDD sky130_fd_sc_hd__fill_2
X_CTS_buf_1_48 _CTS_buf_1_0/A _CTS_buf_1_48/X VSS VDD sky130_fd_sc_hd__clkbuf_4
XANTENNA__1757__A1 _1163_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1518__A _1506_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_77_327 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1253__A SCAN_IN[7] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1693__B1 _1687_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_18_427 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_449 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_235 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_408 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_33_419 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_60_238 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_45_279 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1748__A1 _1152_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1428__A _1430_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1147__B _1139_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0971__A2 _0954_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_7 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_3_22 VSS VDD sky130_fd_sc_hd__fill_2
X_1340_ _1214_/A _1342_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_68_305 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__0986__B _0977_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1271_ _1271_/A SCAN_IN[0] _1274_/A VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_3_88 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_36_202 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_76_382 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1684__B1 _1683_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1922__CLK _1923_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_51_216 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_51_249 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_32_430 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1739__A1 _1144_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0986_ _0953_/X _0977_/X _0982_/X _0986_/D _0986_/X VSS VDD sky130_fd_sc_hd__or4_4
X_1607_ _1601_/X _1607_/B _1608_/B VSS VDD sky130_fd_sc_hd__xor2_4
XANTENNA__1057__B _1057_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__0962__A2 _0961_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_327 VSS VDD sky130_fd_sc_hd__fill_1
X_1538_ _1609_/A _1539_/B VSS VDD sky130_fd_sc_hd__inv_8
X_1469_ _1469_/A _1419_/B _1469_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_67_360 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_408 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1520__B _1520_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1248__A SCAN_IN[9] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1893__D _1893_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_12_97 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0953__A2 _0945_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_5_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_2_367 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_73_352 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1130__A2 _1117_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1666__B1 _1664_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_73_363 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_227 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_430 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_14_441 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_26_290 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1430__B _1422_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_33_249 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1433__A3 _1428_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_41_293 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__0997__A _0996_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_102 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_3 VSS VDD sky130_fd_sc_hd__fill_2
X_1323_ _1894_/Q _1291_/X _1322_/X _1323_/Y VSS VDD sky130_fd_sc_hd__o21ai_4
XANTENNA__1605__B _1605_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1254_ _1155_/A _1579_/B _1254_/X VSS VDD sky130_fd_sc_hd__and2_4
XFILLER_49_371 VSS VDD sky130_fd_sc_hd__decap_8
X_1185_ _1908_/Q _1186_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_24_205 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1404__A1_N _1393_/X VSS VDD sky130_fd_sc_hd__diode_2
X_0969_ _0964_/Y _0959_/Y _0967_/Y _0968_/X _0969_/X VSS VDD sky130_fd_sc_hd__a211o_4
XANTENNA__1188__A2 _1171_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1068__A _1870_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_3_109 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_58_16 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1345__C1 _1344_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_113 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1515__B _1524_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_74_15 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_74_59 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1531__A _1796_/B VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1648__B1 _1602_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_55_341 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1112__A2 _1106_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1888__D _1502_/X VSS VDD sky130_fd_sc_hd__diode_2
XPHY_701 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_355 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_767 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_411 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_282 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1415__A3 _1409_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_404 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1859__RESET_B _1847_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_7_426 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1706__A _1587_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_78_433 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_38_308 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_48_93 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1639__B1 _1580_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_46_341 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_73_160 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_78 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_0_56 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_61_322 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_61_355 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1811__B1 _1796_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1872_ _1173_/X _1872_/Q _1847_/X _1886_/CLK VSS VDD sky130_fd_sc_hd__dfstp_4
XFILLER_9_98 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1319__C _1318_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1590__A2 _1272_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_400 VSS VDD sky130_fd_sc_hd__decap_12
X_1306_ _1276_/A _1305_/X _1276_/A _1305_/X _1306_/Y VSS VDD sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__1351__A SCAN_IN[17] VSS VDD sky130_fd_sc_hd__diode_2
X_1237_ _1237_/A _1241_/A VSS VDD sky130_fd_sc_hd__inv_8
XFILLER_71_119 VSS VDD sky130_fd_sc_hd__decap_3
X_1168_ _1166_/A _1157_/X _1167_/Y _1168_/X VSS VDD sky130_fd_sc_hd__a21o_4
XANTENNA__1645__A3 _1643_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1046__B1_N _1045_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1070__B _1068_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_44_29 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_52_366 VSS VDD sky130_fd_sc_hd__fill_2
X_1099_ _1098_/Y _1245_/A VSS VDD sky130_fd_sc_hd__buf_1
XFILLER_12_219 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1802__B1 _1800_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_20_263 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_274 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_4_429 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_69_48 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_69_15 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1030__A1 _1013_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_79_208 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1245__B _1245_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_75_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_28_330 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_341 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA__1261__A _1127_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_47_149 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_62_119 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_300 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_43_322 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_34_40 VSS VDD sky130_fd_sc_hd__decap_3
XPHY_553 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_285 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_7_245 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1436__A _1384_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_59_70 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_78_296 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_38_105 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_38_127 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_75_91 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1171__A _1170_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_53_108 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_19_352 VSS VDD sky130_fd_sc_hd__fill_2
X_1022_ _1014_/A _1022_/B _1022_/C _1022_/X VSS VDD sky130_fd_sc_hd__and3_4
XANTENNA__1088__A1 _1064_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1088__B2 _1087_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_19_385 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_377 VSS VDD sky130_fd_sc_hd__decap_12
X_1924_ _1846_/Y _1924_/Q RESET_N _1924_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
XANTENNA__1260__A1 _1430_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1855_ _1855_/D _0955_/A _1847_/X _1853_/CLK VSS VDD sky130_fd_sc_hd__dfrtp_4
X_1786_ _1620_/X _1786_/B _1786_/Y VSS VDD sky130_fd_sc_hd__nor2_4
XANTENNA__1049__C _1048_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1346__A SCAN_IN[20] VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1563__A2 _1796_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_241 VSS VDD sky130_fd_sc_hd__decap_3
XANTENNA__1315__A2 _1314_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_69_296 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_57_425 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1079__A1 _1874_/Q VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1512__C _1510_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1081__A _1081_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1079__B2 _0991_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_25_355 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_40_369 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_4_215 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1003__A1 _0963_/Y VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1554__A2 _1613_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1256__A _1255_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_4_259 VSS VDD sky130_fd_sc_hd__decap_12
XFILLER_20_53 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_20_64 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_0_443 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_29_62 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1703__B _1703_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_48_447 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_63_428 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_300 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_182 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1490__A1 _1461_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1490__B2 _1489_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_303 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_43_174 VSS VDD sky130_fd_sc_hd__fill_2
XPHY_350 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VSS VDD sky130_fd_sc_hd__decap_4
XPHY_372 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1793__A2 _1743_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1640_ _1734_/A _1634_/X _1640_/X VSS VDD sky130_fd_sc_hd__or2_4
XFILLER_6_11 VSS VDD sky130_fd_sc_hd__decap_3
X_1571_ _1571_/A _1571_/B _1571_/X VSS VDD sky130_fd_sc_hd__or2_4
XANTENNA__1166__A _1166_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_6_88 VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_3 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_39_425 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_66_255 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_160 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_19_171 VSS VDD sky130_fd_sc_hd__decap_12
X_1005_ _1005_/A _1005_/Y VSS VDD sky130_fd_sc_hd__inv_8
XANTENNA__1481__A1 _1304_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1481__B2 _1480_/X VSS VDD sky130_fd_sc_hd__diode_2
X_1907_ _1907_/D _1772_/A _1847_/X _1924_/Q VSS VDD sky130_fd_sc_hd__dfstp_4
XANTENNA__1233__B2 _1451_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1784__A2 _1759_/A VSS VDD sky130_fd_sc_hd__diode_2
X_1838_ _1837_/A _1836_/C _1839_/C VSS VDD sky130_fd_sc_hd__nand2_4
X_1769_ _1769_/A _1716_/B _1716_/C _1769_/Y VSS VDD sky130_fd_sc_hd__nor3_4
XANTENNA__1076__A _1873_/Q VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_1_229 VSS VDD sky130_fd_sc_hd__fill_1
XANTENNA__1804__A _1803_/C VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_66_49 VSS VDD sky130_fd_sc_hd__decap_6
XANTENNA__1523__B _1523_/B VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_57_288 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_45_428 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_72_247 VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_141 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_15_20 VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_163 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_13_336 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_15_75 VSS VDD sky130_fd_sc_hd__decap_8
XANTENNA__1896__D _1896_/D VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_15_97 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_21_380 VSS VDD sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_0_16_A _CTS_buf_1_16/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1224__B2 _1215_/A VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1775__A2 _1769_/Y VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_31_74 VSS VDD sky130_fd_sc_hd__decap_4
XANTENNA__1527__A2 _1492_/X VSS VDD sky130_fd_sc_hd__diode_2
XANTENNA__1714__A _1689_/A VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_0_273 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_63_225 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_93 VSS VDD sky130_fd_sc_hd__fill_2
XFILLER_56_82 VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_152 VSS VDD sky130_fd_sc_hd__fill_1
XFILLER_16_163 VSS VDD sky130_fd_sc_hd__decap_8
XPHY_180 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1766__A2 _1696_/X VSS VDD sky130_fd_sc_hd__diode_2
XFILLER_68_3 VSS VDD sky130_fd_sc_hd__fill_2
XANTENNA__1608__B _1608_/B VSS VDD sky130_fd_sc_hd__diode_2
X_1623_ _1694_/A _1618_/Y _1591_/X _1622_/Y _1623_/X VSS VDD sky130_fd_sc_hd__a211o_4
XANTENNA__1851__CLK _1865_/CLK VSS VDD sky130_fd_sc_hd__diode_2
X_1554_ _1131_/X _1613_/A _1551_/X _1553_/X _1554_/X VSS VDD sky130_fd_sc_hd__o22a_4
X_1485_ _1430_/A _1427_/A _1478_/X _1484_/X _1485_/Y VSS VDD sky130_fd_sc_hd__a22oi_4
.ends

