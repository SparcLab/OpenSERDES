VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

MACRO CLK_RECOVERY
  CLASS BLOCK ;
  FOREIGN CLK_RECOVERY ;
  ORIGIN 0.000 0.000 ;
  SIZE 228.850 BY 239.570 ;
  PIN BB_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 235.570 40.850 239.570 ;
    END
  END BB_IN
  PIN CLK_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END CLK_IN
  PIN CLK_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END CLK_OUT
  PIN DATA_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END DATA_OUT
  PIN RESET_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.070 235.570 98.350 239.570 ;
    END
  END RESET_N
  PIN SCAN_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 46.960 228.850 47.560 ;
    END
  END SCAN_IN[0]
  PIN SCAN_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 131.960 228.850 132.560 ;
    END
  END SCAN_IN[10]
  PIN SCAN_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END SCAN_IN[11]
  PIN SCAN_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END SCAN_IN[12]
  PIN SCAN_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.990 235.570 214.270 239.570 ;
    END
  END SCAN_IN[13]
  PIN SCAN_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END SCAN_IN[14]
  PIN SCAN_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 235.570 11.870 239.570 ;
    END
  END SCAN_IN[15]
  PIN SCAN_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 174.800 228.850 175.400 ;
    END
  END SCAN_IN[16]
  PIN SCAN_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 89.120 228.850 89.720 ;
    END
  END SCAN_IN[17]
  PIN SCAN_IN[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END SCAN_IN[18]
  PIN SCAN_IN[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END SCAN_IN[19]
  PIN SCAN_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 235.570 127.330 239.570 ;
    END
  END SCAN_IN[1]
  PIN SCAN_IN[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END SCAN_IN[20]
  PIN SCAN_IN[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 235.570 69.830 239.570 ;
    END
  END SCAN_IN[21]
  PIN SCAN_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END SCAN_IN[2]
  PIN SCAN_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.030 235.570 156.310 239.570 ;
    END
  END SCAN_IN[3]
  PIN SCAN_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 4.120 228.850 4.720 ;
    END
  END SCAN_IN[4]
  PIN SCAN_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END SCAN_IN[5]
  PIN SCAN_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.010 235.570 185.290 239.570 ;
    END
  END SCAN_IN[6]
  PIN SCAN_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END SCAN_IN[7]
  PIN SCAN_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END SCAN_IN[8]
  PIN SCAN_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 224.850 217.640 228.850 218.240 ;
    END
  END SCAN_IN[9]
  PIN VDD
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 223.100 28.090 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 223.100 104.680 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 223.100 228.565 ;
      LAYER met1 ;
        RECT 0.070 0.380 223.100 235.580 ;
      LAYER met2 ;
        RECT 5.610 235.290 11.310 235.690 ;
        RECT 12.150 235.290 40.290 235.690 ;
        RECT 41.130 235.290 69.270 235.690 ;
        RECT 70.110 235.290 97.790 235.690 ;
        RECT 98.630 235.290 126.770 235.690 ;
        RECT 127.610 235.290 155.750 235.690 ;
        RECT 156.590 235.290 184.730 235.690 ;
        RECT 185.570 235.290 213.710 235.690 ;
        RECT 214.550 235.290 224.390 235.690 ;
        RECT 5.610 4.280 224.390 235.290 ;
        RECT 5.610 0.270 28.330 4.280 ;
        RECT 29.170 0.270 57.310 4.280 ;
        RECT 58.150 0.270 86.290 4.280 ;
        RECT 87.130 0.270 115.270 4.280 ;
        RECT 116.110 0.270 144.250 4.280 ;
        RECT 145.090 0.270 173.230 4.280 ;
        RECT 174.070 0.270 202.210 4.280 ;
        RECT 203.050 0.270 224.390 4.280 ;
      LAYER met3 ;
        RECT 0.270 218.640 224.850 228.645 ;
        RECT 0.270 217.240 224.450 218.640 ;
        RECT 0.270 214.560 224.850 217.240 ;
        RECT 4.400 213.160 224.850 214.560 ;
        RECT 0.270 175.800 224.850 213.160 ;
        RECT 0.270 174.400 224.450 175.800 ;
        RECT 0.270 171.720 224.850 174.400 ;
        RECT 4.400 170.320 224.850 171.720 ;
        RECT 0.270 132.960 224.850 170.320 ;
        RECT 0.270 131.560 224.450 132.960 ;
        RECT 0.270 128.880 224.850 131.560 ;
        RECT 4.400 127.480 224.850 128.880 ;
        RECT 0.270 90.120 224.850 127.480 ;
        RECT 0.270 88.720 224.450 90.120 ;
        RECT 0.270 86.040 224.850 88.720 ;
        RECT 4.400 84.640 224.850 86.040 ;
        RECT 0.270 47.960 224.850 84.640 ;
        RECT 0.270 46.560 224.450 47.960 ;
        RECT 0.270 43.200 224.850 46.560 ;
        RECT 4.400 41.800 224.850 43.200 ;
        RECT 0.270 5.120 224.850 41.800 ;
        RECT 0.270 4.255 224.450 5.120 ;
      LAYER met4 ;
        RECT 0.295 10.640 176.240 228.720 ;
      LAYER met5 ;
        RECT 5.520 179.670 223.100 181.270 ;
  END
END CLK_RECOVERY
END LIBRARY

