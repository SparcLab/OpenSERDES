/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */
/* With case-insensitive names (SPICE-compatible) */

module serializer_unit_cell_1(
    inout vpwr,
    inout vgnd,
    input CLK,
    output COMPLETE,
    output INTERNAL_FINISH,
    input READY,
    input RESET,
    output SERIAL_OUT,
    input VDD,
    input VSS,
    output [5:0] COUNT,
    input [31:0] PAR_IN1,
    input [31:0] PAR_IN2,
    input [31:0] PAR_IN3,
    input [31:0] PAR_IN4,
    input [31:0] PAR_IN5,
    input [31:0] PAR_IN6,
    input [31:0] PAR_IN7,
    input [31:0] PAR_IN8,
    output [3:0] SAMPLE_COUNT
);

wire _0472_ ;
wire _0052_ ;
wire _0108_ ;
wire _0281_ ;
wire _0337_ ;
wire _0090_ ;
wire _0146_ ;
wire _0375_ ;
wire _0184_ ;
wire _0469_ ;
wire _0049_ ;
wire _0278_ ;
wire _0087_ ;
wire _0202_ ;
wire _0431_ ;
wire _0011_ ;
wire _0240_ ;
wire _0105_ ;
wire _0334_ ;
wire _0143_ ;
wire _0372_ ;
wire _0428_ ;
wire _0008_ ;
wire _0181_ ;
wire _0237_ ;
wire _0466_ ;
wire _0046_ ;
wire _0275_ ;
wire _0084_ ;
wire _0369_ ;
wire _0178_ ;
wire READY ;
wire [3:0] SAMPLE_COUNT ;
wire _0102_ ;
wire SERIAL_OUT ;
wire _0331_ ;
wire _0140_ ;
wire _0425_ ;
wire _0005_ ;
wire _0234_ ;
wire _0463_ ;
wire _0043_ ;
wire _0272_ ;
wire _0328_ ;
wire _0081_ ;
wire _0137_ ;
wire _0366_ ;
wire _0175_ ;
wire _0269_ ;
wire _0498_ ;
wire _0078_ ;
wire _0422_ ;
wire _0002_ ;
wire _0231_ ;
wire _0460_ ;
wire _0040_ ;
wire _0325_ ;
wire _0134_ ;
wire _0363_ ;
wire _0419_ ;
wire _0172_ ;
wire _0228_ ;
wire _0457_ ;
wire _0037_ ;
wire _0266_ ;
wire _0495_ ;
wire _0075_ ;
wire _0169_ ;
wire _0398_ ;
wire RESET ;
wire _0322_ ;
wire _0131_ ;
wire _0360_ ;
wire _0416_ ;
wire _0225_ ;
wire _0454_ ;
wire _0034_ ;
wire _0263_ ;
wire _0319_ ;
wire _0492_ ;
wire _0072_ ;
wire _0128_ ;
wire _0357_ ;
wire _0166_ ;
wire _0395_ ;
wire _0489_ ;
wire _0069_ ;
wire _0298_ ;
wire _0413_ ;
wire _0222_ ;
wire _0451_ ;
wire _0031_ ;
wire _0507_ ;
wire _0260_ ;
wire _0316_ ;
wire _0125_ ;
wire _0354_ ;
wire _0163_ ;
wire _0219_ ;
wire _0392_ ;
wire _0448_ ;
wire _0028_ ;
wire _0257_ ;
wire _0486_ ;
wire _0066_ ;
wire _0295_ ;
wire _0389_ ;
wire _0198_ ;
wire _0410_ ;
wire _0504_ ;
wire _0313_ ;
wire _0122_ ;
wire _0351_ ;
wire clknet_1_1_0_CLK ;
wire _0407_ ;
wire _0160_ ;
wire _0216_ ;
wire _0445_ ;
wire _0025_ ;
wire _0254_ ;
wire _0483_ ;
wire _0063_ ;
wire _0119_ ;
wire _0292_ ;
wire _0348_ ;
wire _0157_ ;
wire _0386_ ;
wire VSS ;
wire _0195_ ;
wire _0289_ ;
wire _0501_ ;
wire _0098_ ;
wire _0310_ ;
wire _0404_ ;
wire _0213_ ;
wire _0442_ ;
wire _0022_ ;
wire _0251_ ;
wire _0307_ ;
wire _0480_ ;
wire _0060_ ;
wire _0116_ ;
wire _0345_ ;
wire _0154_ ;
wire _0383_ ;
wire _0439_ ;
wire _0019_ ;
wire _0192_ ;
wire _0248_ ;
wire _0477_ ;
wire _0057_ ;
wire _0286_ ;
wire _0095_ ;
wire _0189_ ;
wire _0401_ ;
wire _0210_ ;
wire _0304_ ;
wire _0113_ ;
wire _0342_ ;
wire _0151_ ;
wire _0207_ ;
wire _0380_ ;
wire _0436_ ;
wire _0016_ ;
wire _0245_ ;
wire _0474_ ;
wire _0054_ ;
wire _0283_ ;
wire _0339_ ;
wire _0092_ ;
wire _0148_ ;
wire _0377_ ;
wire _0186_ ;
wire _0089_ ;
wire _0301_ ;
wire _0110_ ;
wire _0204_ ;
wire _0433_ ;
wire _0013_ ;
wire _0242_ ;
wire _0471_ ;
wire _0051_ ;
wire _0107_ ;
wire _0280_ ;
wire _0336_ ;
wire _0145_ ;
wire _0374_ ;
wire _0183_ ;
wire _0239_ ;
wire _0468_ ;
wire _0048_ ;
wire _0277_ ;
wire _0086_ ;
wire _0201_ ;
wire _0430_ ;
wire _0010_ ;
wire _0104_ ;
wire _0333_ ;
wire _0142_ ;
wire _0371_ ;
wire _0427_ ;
wire _0007_ ;
wire _0180_ ;
wire _0236_ ;
wire _0465_ ;
wire _0045_ ;
wire _0274_ ;
wire _0083_ ;
wire _0139_ ;
wire _0368_ ;
wire _0177_ ;
wire VDD ;
wire _0101_ ;
wire _0330_ ;
wire _0424_ ;
wire _0004_ ;
wire _0233_ ;
wire _0462_ ;
wire _0042_ ;
wire _0271_ ;
wire _0327_ ;
wire _0080_ ;
wire _0136_ ;
wire _0365_ ;
wire _0174_ ;
wire _0459_ ;
wire _0039_ ;
wire _0268_ ;
wire _0497_ ;
wire _0077_ ;
wire _0421_ ;
wire _0001_ ;
wire _0230_ ;
wire _0324_ ;
wire _0133_ ;
wire _0362_ ;
wire _0418_ ;
wire _0171_ ;
wire _0227_ ;
wire _0456_ ;
wire _0036_ ;
wire _0265_ ;
wire _0494_ ;
wire _0074_ ;
wire _0359_ ;
wire _0168_ ;
wire _0397_ ;
wire _0321_ ;
wire _0130_ ;
wire _0415_ ;
wire _0224_ ;
wire _0453_ ;
wire _0033_ ;
wire _0262_ ;
wire _0318_ ;
wire _0491_ ;
wire _0071_ ;
wire _0127_ ;
wire _0356_ ;
wire _0165_ ;
wire _0394_ ;
wire _0259_ ;
wire _0488_ ;
wire _0068_ ;
wire _0297_ ;
wire _0412_ ;
wire _0221_ ;
wire _0450_ ;
wire _0030_ ;
wire _0506_ ;
wire _0315_ ;
wire _0124_ ;
wire _0353_ ;
wire _0409_ ;
wire _0162_ ;
wire _0218_ ;
wire _0391_ ;
wire _0447_ ;
wire _0027_ ;
wire _0256_ ;
wire _0485_ ;
wire _0065_ ;
wire _0294_ ;
wire _0159_ ;
wire _0388_ ;
wire _0197_ ;
wire _0503_ ;
wire _0312_ ;
wire _0121_ ;
wire _0350_ ;
wire _0406_ ;
wire _0215_ ;
wire _0444_ ;
wire _0024_ ;
wire _0253_ ;
wire _0309_ ;
wire _0482_ ;
wire _0062_ ;
wire _0118_ ;
wire _0291_ ;
wire _0347_ ;
wire _0156_ ;
wire _0385_ ;
wire _0194_ ;
wire _0479_ ;
wire _0059_ ;
wire _0288_ ;
wire _0500_ ;
wire _0097_ ;
wire _0403_ ;
wire _0212_ ;
wire _0441_ ;
wire _0021_ ;
wire _0250_ ;
wire _0306_ ;
wire _0115_ ;
wire _0344_ ;
wire _0153_ ;
wire _0209_ ;
wire _0382_ ;
wire _0438_ ;
wire _0018_ ;
wire _0191_ ;
wire _0247_ ;
wire INTERNAL_FINISH ;
wire _0476_ ;
wire _0056_ ;
wire _0285_ ;
wire _0094_ ;
wire _0379_ ;
wire _0188_ ;
wire _0400_ ;
wire _0303_ ;
wire _0112_ ;
wire _0341_ ;
wire [31:0] PAR_IN1 ;
wire [31:0] PAR_IN2 ;
wire [31:0] PAR_IN3 ;
wire [31:0] PAR_IN4 ;
wire [31:0] PAR_IN5 ;
wire [31:0] PAR_IN6 ;
wire [31:0] PAR_IN7 ;
wire [31:0] PAR_IN8 ;
wire _0150_ ;
wire _0206_ ;
wire CLK ;
wire _0435_ ;
wire _0015_ ;
wire _0244_ ;
wire _0473_ ;
wire _0053_ ;
wire _0109_ ;
wire _0282_ ;
wire _0338_ ;
wire _0091_ ;
wire _0147_ ;
wire _0376_ ;
wire _0185_ ;
wire _0279_ ;
wire _0088_ ;
wire _0300_ ;
wire _0203_ ;
wire _0432_ ;
wire _0012_ ;
wire _0241_ ;
wire _0470_ ;
wire _0050_ ;
wire _0106_ ;
wire _0335_ ;
wire _0144_ ;
wire _0373_ ;
wire _0429_ ;
wire _0009_ ;
wire _0182_ ;
wire _0238_ ;
wire _0467_ ;
wire _0047_ ;
wire _0276_ ;
wire _0085_ ;
wire _0179_ ;
wire _0200_ ;
wire _0103_ ;
wire _0332_ ;
wire _0141_ ;
wire _0370_ ;
wire _0426_ ;
wire _0006_ ;
wire _0235_ ;
wire _0464_ ;
wire _0044_ ;
wire _0273_ ;
wire _0329_ ;
wire _0082_ ;
wire _0138_ ;
wire _0367_ ;
wire _0176_ ;
wire _0499_ ;
wire _0079_ ;
wire _0100_ ;
wire clknet_1_0_0_CLK ;
wire _0423_ ;
wire _0003_ ;
wire _0232_ ;
wire _0461_ ;
wire _0041_ ;
wire clknet_0_CLK ;
wire _0270_ ;
wire _0326_ ;
wire _0135_ ;
wire _0364_ ;
wire _0173_ ;
wire _0229_ ;
wire _0458_ ;
wire _0038_ ;
wire _0267_ ;
wire _0496_ ;
wire _0076_ ;
wire _0399_ ;
wire COMPLETE ;
wire _0420_ ;
wire _0000_ ;
wire _0323_ ;
wire _0132_ ;
wire _0361_ ;
wire _0417_ ;
wire _0170_ ;
wire _0226_ ;
wire _0455_ ;
wire _0035_ ;
wire _0264_ ;
wire _0493_ ;
wire _0073_ ;
wire _0129_ ;
wire [5:0] COUNT ;
wire _0358_ ;
wire _0167_ ;
wire _0396_ ;
wire _0299_ ;
wire _0320_ ;
wire _0414_ ;
wire _0223_ ;
wire _0452_ ;
wire _0032_ ;
wire _0261_ ;
wire _0317_ ;
wire _0490_ ;
wire _0070_ ;
wire _0126_ ;
wire _0355_ ;
wire _0164_ ;
wire _0393_ ;
wire _0449_ ;
wire _0029_ ;
wire _0258_ ;
wire _0487_ ;
wire _0067_ ;
wire _0296_ ;
wire _0199_ ;
wire _0411_ ;
wire _0220_ ;
wire _0505_ ;
wire _0314_ ;
wire _0123_ ;
wire _0352_ ;
wire _0408_ ;
wire _0161_ ;
wire _0217_ ;
wire _0390_ ;
wire _0446_ ;
wire _0026_ ;
wire _0255_ ;
wire _0484_ ;
wire _0064_ ;
wire _0293_ ;
wire _0349_ ;
wire _0158_ ;
wire _0387_ ;
wire _0196_ ;
wire _0502_ ;
wire _0099_ ;
wire _0311_ ;
wire _0120_ ;
wire _0405_ ;
wire _0214_ ;
wire _0443_ ;
wire _0023_ ;
wire _0252_ ;
wire _0308_ ;
wire _0481_ ;
wire _0061_ ;
wire _0117_ ;
wire _0290_ ;
wire _0346_ ;
wire _0155_ ;
wire _0384_ ;
wire _0193_ ;
wire _0249_ ;
wire _0478_ ;
wire _0058_ ;
wire _0287_ ;
wire _0096_ ;
wire _0402_ ;
wire _0211_ ;
wire _0440_ ;
wire _0020_ ;
wire _0305_ ;
wire _0114_ ;
wire _0343_ ;
wire _0152_ ;
wire _0208_ ;
wire _0381_ ;
wire _0437_ ;
wire _0017_ ;
wire _0190_ ;
wire _0246_ ;
wire _0475_ ;
wire _0055_ ;
wire _0284_ ;
wire _0093_ ;
wire _0149_ ;
wire _0378_ ;
wire _0187_ ;
wire _0302_ ;
wire _0111_ ;
wire _0340_ ;
wire _0205_ ;
wire _0434_ ;
wire _0014_ ;
wire _0243_ ;

sky130_fd_sc_hd__buf_1 _0508_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[0]),
    .X(_0013_)
);

sky130_fd_sc_hd__inv_8 _0509_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[4]),
    .Y(_0014_)
);

sky130_fd_sc_hd__buf_1 _0510_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0014_),
    .X(_0015_)
);

sky130_fd_sc_hd__buf_1 _0511_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0015_),
    .X(_0016_)
);

sky130_fd_sc_hd__buf_1 _0512_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0016_),
    .X(_0017_)
);

sky130_fd_sc_hd__inv_8 _0513_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[3]),
    .Y(_0018_)
);

sky130_fd_sc_hd__buf_1 _0514_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0018_),
    .X(_0019_)
);

sky130_fd_sc_hd__inv_8 _0515_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[2]),
    .Y(_0020_)
);

sky130_fd_sc_hd__inv_8 _0516_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[0]),
    .Y(_0021_)
);

sky130_fd_sc_hd__inv_8 _0517_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[1]),
    .Y(_0022_)
);

sky130_fd_sc_hd__or2_4 _0518_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0021_),
    .B(_0022_),
    .X(_0023_)
);

sky130_fd_sc_hd__or2_4 _0519_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0020_),
    .B(_0023_),
    .X(_0024_)
);

sky130_fd_sc_hd__or2_4 _0520_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0019_),
    .B(_0024_),
    .X(_0025_)
);

sky130_fd_sc_hd__inv_8 _0521_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[5]),
    .Y(_0026_)
);

sky130_fd_sc_hd__o21a_4 _0522_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0017_),
    .A2(_0025_),
    .B1(_0026_),
    .X(_0027_)
);

sky130_fd_sc_hd__buf_1 _0523_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0027_),
    .X(_0028_)
);

sky130_fd_sc_hd__inv_8 _0524_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0028_),
    .Y(_0029_)
);

sky130_fd_sc_hd__inv_8 _0525_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[3]),
    .Y(_0030_)
);

sky130_fd_sc_hd__buf_1 _0526_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0030_),
    .X(_0031_)
);

sky130_fd_sc_hd__buf_1 _0527_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0031_),
    .X(_0032_)
);

sky130_fd_sc_hd__inv_8 _0528_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COMPLETE),
    .Y(_0033_)
);

sky130_fd_sc_hd__buf_1 _0529_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0033_),
    .X(_0034_)
);

sky130_fd_sc_hd__and4_4 _0530_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0013_),
    .B(_0029_),
    .C(_0032_),
    .D(_0034_),
    .X(_0035_)
);

sky130_fd_sc_hd__inv_8 _0531_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(INTERNAL_FINISH),
    .Y(_0036_)
);

sky130_fd_sc_hd__o21a_4 _0532_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0032_),
    .A2(_0036_),
    .B1(READY),
    .X(_0037_)
);

sky130_fd_sc_hd__inv_8 _0533_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0037_),
    .Y(_0038_)
);

sky130_fd_sc_hd__buf_1 _0534_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0038_),
    .X(_0039_)
);

sky130_fd_sc_hd__buf_1 _0535_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COMPLETE),
    .X(_0040_)
);

sky130_fd_sc_hd__and2_4 _0536_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0032_),
    .B(_0028_),
    .X(_0041_)
);

sky130_fd_sc_hd__inv_8 _0537_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[0]),
    .Y(_0042_)
);

sky130_fd_sc_hd__buf_1 _0538_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0042_),
    .X(_0043_)
);

sky130_fd_sc_hd__o21a_4 _0539_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0040_),
    .A2(_0041_),
    .B1(_0043_),
    .X(_0044_)
);

sky130_fd_sc_hd__nor3_4 _0540_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0035_),
    .B(_0039_),
    .C(_0044_),
    .Y(_0008_)
);

sky130_fd_sc_hd__buf_1 _0541_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[3]),
    .X(_0045_)
);

sky130_fd_sc_hd__buf_1 _0542_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[1]),
    .X(_0046_)
);

sky130_fd_sc_hd__and3_4 _0543_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0046_),
    .B(_0013_),
    .C(_0029_),
    .X(_0047_)
);

sky130_fd_sc_hd__inv_8 _0544_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[1]),
    .Y(_0048_)
);

sky130_fd_sc_hd__buf_1 _0545_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0048_),
    .X(_0049_)
);

sky130_fd_sc_hd__o21a_4 _0546_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0043_),
    .A2(_0028_),
    .B1(_0049_),
    .X(_0050_)
);

sky130_fd_sc_hd__or3_4 _0547_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0045_),
    .B(_0047_),
    .C(_0050_),
    .X(_0051_)
);

sky130_fd_sc_hd__a21o_4 _0548_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0049_),
    .A2(_0040_),
    .B1(_0039_),
    .X(_0052_)
);

sky130_fd_sc_hd__a21oi_4 _0549_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0034_),
    .A2(_0051_),
    .B1(_0052_),
    .Y(_0009_)
);

sky130_fd_sc_hd__buf_1 _0550_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0045_),
    .X(_0053_)
);

sky130_fd_sc_hd__buf_1 _0551_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[2]),
    .X(_0054_)
);

sky130_fd_sc_hd__and2_4 _0552_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0033_),
    .B(_0047_),
    .X(_0055_)
);

sky130_fd_sc_hd__nor2_4 _0553_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0054_),
    .B(_0055_),
    .Y(_0056_)
);

sky130_fd_sc_hd__and2_4 _0554_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0054_),
    .B(_0055_),
    .X(_0057_)
);

sky130_fd_sc_hd__a2111oi_4 _0555_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0053_),
    .A2(_0034_),
    .B1(_0039_),
    .C1(_0056_),
    .D1(_0057_),
    .Y(_0010_)
);

sky130_fd_sc_hd__o21a_4 _0556_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0053_),
    .A2(_0057_),
    .B1(_0037_),
    .X(_0011_)
);

sky130_fd_sc_hd__o21a_4 _0557_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0045_),
    .A2(COUNT[5]),
    .B1(_0021_),
    .X(_0058_)
);

sky130_fd_sc_hd__a2111oi_4 _0558_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0032_),
    .A2(COUNT[0]),
    .B1(_0058_),
    .C1(_0040_),
    .D1(_0039_),
    .Y(_0001_)
);

sky130_fd_sc_hd__buf_1 _0559_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0032_),
    .X(_0059_)
);

sky130_fd_sc_hd__o21a_4 _0560_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(COUNT[0]),
    .A2(COUNT[1]),
    .B1(_0023_),
    .X(_0060_)
);

sky130_fd_sc_hd__nand2_4 _0561_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0028_),
    .B(_0060_),
    .Y(_0061_)
);

sky130_fd_sc_hd__or2_4 _0562_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COMPLETE),
    .B(_0038_),
    .X(_0062_)
);

sky130_fd_sc_hd__a21o_4 _0563_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0053_),
    .A2(_0022_),
    .B1(_0062_),
    .X(_0063_)
);

sky130_fd_sc_hd__a21oi_4 _0564_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0059_),
    .A2(_0061_),
    .B1(_0063_),
    .Y(_0002_)
);

sky130_fd_sc_hd__buf_1 _0565_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0020_),
    .X(_0064_)
);

sky130_fd_sc_hd__inv_8 _0566_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0024_),
    .Y(_0065_)
);

sky130_fd_sc_hd__a211o_4 _0567_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0064_),
    .A2(_0023_),
    .B1(_0065_),
    .C1(_0029_),
    .X(_0066_)
);

sky130_fd_sc_hd__a21o_4 _0568_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0053_),
    .A2(_0064_),
    .B1(_0062_),
    .X(_0067_)
);

sky130_fd_sc_hd__a21oi_4 _0569_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0059_),
    .A2(_0066_),
    .B1(_0067_),
    .Y(_0003_)
);

sky130_fd_sc_hd__buf_1 _0570_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[3]),
    .X(_0068_)
);

sky130_fd_sc_hd__buf_1 _0571_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0068_),
    .X(_0069_)
);

sky130_fd_sc_hd__o21a_4 _0572_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0069_),
    .A2(_0065_),
    .B1(_0025_),
    .X(_0070_)
);

sky130_fd_sc_hd__nand2_4 _0573_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0028_),
    .B(_0070_),
    .Y(_0071_)
);

sky130_fd_sc_hd__buf_1 _0574_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0019_),
    .X(_0072_)
);

sky130_fd_sc_hd__a21o_4 _0575_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0045_),
    .A2(_0072_),
    .B1(_0062_),
    .X(_0073_)
);

sky130_fd_sc_hd__a21oi_4 _0576_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0059_),
    .A2(_0071_),
    .B1(_0073_),
    .Y(_0004_)
);

sky130_fd_sc_hd__or2_4 _0577_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0045_),
    .B(_0025_),
    .X(_0074_)
);

sky130_fd_sc_hd__a21o_4 _0578_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0017_),
    .A2(_0074_),
    .B1(_0062_),
    .X(_0075_)
);

sky130_fd_sc_hd__a21oi_4 _0579_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0059_),
    .A2(_0029_),
    .B1(_0075_),
    .Y(_0005_)
);

sky130_fd_sc_hd__and4_4 _0580_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0053_),
    .B(_0034_),
    .C(COUNT[5]),
    .D(_0037_),
    .X(_0006_)
);

sky130_fd_sc_hd__and4_4 _0581_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0059_),
    .B(_0054_),
    .C(READY),
    .D(_0055_),
    .X(_0000_)
);

sky130_fd_sc_hd__o22a_4 _0582_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0040_),
    .A2(_0041_),
    .B1(_0034_),
    .B2(_0036_),
    .X(_0076_)
);

sky130_fd_sc_hd__nor2_4 _0583_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0039_),
    .B(_0076_),
    .Y(_0007_)
);

sky130_fd_sc_hd__buf_1 _0584_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0015_),
    .X(_0077_)
);

sky130_fd_sc_hd__inv_8 _0585_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[2]),
    .Y(_0078_)
);

sky130_fd_sc_hd__and3_4 _0586_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0048_),
    .B(_0042_),
    .C(_0078_),
    .X(_0079_)
);

sky130_fd_sc_hd__or2_4 _0587_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[3]),
    .B(_0079_),
    .X(_0080_)
);

sky130_fd_sc_hd__buf_1 _0588_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0080_),
    .X(_0081_)
);

sky130_fd_sc_hd__buf_1 _0589_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0081_),
    .X(_0082_)
);

sky130_fd_sc_hd__inv_8 _0590_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0082_),
    .Y(_0083_)
);

sky130_fd_sc_hd__buf_1 _0591_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0083_),
    .X(_0084_)
);

sky130_fd_sc_hd__buf_1 _0592_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0084_),
    .X(_0085_)
);

sky130_fd_sc_hd__or2_4 _0593_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[15]),
    .B(_0085_),
    .X(_0086_)
);

sky130_fd_sc_hd__and4_4 _0594_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0030_),
    .B(SAMPLE_COUNT[2]),
    .C(_0049_),
    .D(_0013_),
    .X(_0087_)
);

sky130_fd_sc_hd__buf_1 _0595_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0087_),
    .X(_0088_)
);

sky130_fd_sc_hd__buf_1 _0596_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0088_),
    .X(_0089_)
);

sky130_fd_sc_hd__buf_1 _0597_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0089_),
    .X(_0090_)
);

sky130_fd_sc_hd__and4_4 _0598_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0046_),
    .B(SAMPLE_COUNT[0]),
    .C(_0030_),
    .D(_0078_),
    .X(_0091_)
);

sky130_fd_sc_hd__buf_1 _0599_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0091_),
    .X(_0092_)
);

sky130_fd_sc_hd__buf_1 _0600_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0092_),
    .X(_0093_)
);

sky130_fd_sc_hd__and2_4 _0601_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[15]),
    .B(_0093_),
    .X(_0094_)
);

sky130_fd_sc_hd__a21o_4 _0602_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[15]),
    .A2(_0090_),
    .B1(_0094_),
    .X(_0095_)
);

sky130_fd_sc_hd__and4_4 _0603_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0046_),
    .B(_0013_),
    .C(_0030_),
    .D(SAMPLE_COUNT[2]),
    .X(_0096_)
);

sky130_fd_sc_hd__buf_1 _0604_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0096_),
    .X(_0097_)
);

sky130_fd_sc_hd__buf_1 _0605_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0097_),
    .X(_0098_)
);

sky130_fd_sc_hd__buf_1 _0606_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0098_),
    .X(_0099_)
);

sky130_fd_sc_hd__and4_4 _0607_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0031_),
    .B(_0054_),
    .C(_0049_),
    .D(_0043_),
    .X(_0100_)
);

sky130_fd_sc_hd__buf_1 _0608_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0100_),
    .X(_0101_)
);

sky130_fd_sc_hd__buf_1 _0609_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0101_),
    .X(_0102_)
);

sky130_fd_sc_hd__and2_4 _0610_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[15]),
    .B(_0102_),
    .X(_0103_)
);

sky130_fd_sc_hd__a21o_4 _0611_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[15]),
    .A2(_0099_),
    .B1(_0103_),
    .X(_0104_)
);

sky130_fd_sc_hd__and4_4 _0612_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0031_),
    .B(_0078_),
    .C(_0046_),
    .D(_0043_),
    .X(_0105_)
);

sky130_fd_sc_hd__buf_1 _0613_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0105_),
    .X(_0106_)
);

sky130_fd_sc_hd__buf_1 _0614_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0106_),
    .X(_0107_)
);

sky130_fd_sc_hd__buf_1 _0615_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0081_),
    .X(_0108_)
);

sky130_fd_sc_hd__buf_1 _0616_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0108_),
    .X(_0109_)
);

sky130_fd_sc_hd__a21o_4 _0617_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[15]),
    .A2(_0107_),
    .B1(_0109_),
    .X(_0110_)
);

sky130_fd_sc_hd__and4_4 _0618_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0031_),
    .B(_0078_),
    .C(_0049_),
    .D(_0013_),
    .X(_0111_)
);

sky130_fd_sc_hd__buf_1 _0619_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0111_),
    .X(_0112_)
);

sky130_fd_sc_hd__buf_1 _0620_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0112_),
    .X(_0113_)
);

sky130_fd_sc_hd__and4_4 _0621_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0031_),
    .B(_0054_),
    .C(_0046_),
    .D(_0043_),
    .X(_0114_)
);

sky130_fd_sc_hd__buf_1 _0622_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0114_),
    .X(_0115_)
);

sky130_fd_sc_hd__buf_1 _0623_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0115_),
    .X(_0116_)
);

sky130_fd_sc_hd__and2_4 _0624_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[15]),
    .B(_0116_),
    .X(_0117_)
);

sky130_fd_sc_hd__a21o_4 _0625_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[15]),
    .A2(_0113_),
    .B1(_0117_),
    .X(_0118_)
);

sky130_fd_sc_hd__or4_4 _0626_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0095_),
    .B(_0104_),
    .C(_0110_),
    .D(_0118_),
    .X(_0119_)
);

sky130_fd_sc_hd__and3_4 _0627_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0077_),
    .B(_0086_),
    .C(_0119_),
    .X(_0120_)
);

sky130_fd_sc_hd__buf_1 _0628_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[4]),
    .X(_0121_)
);

sky130_fd_sc_hd__buf_1 _0629_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0121_),
    .X(_0122_)
);

sky130_fd_sc_hd__buf_1 _0630_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0084_),
    .X(_0123_)
);

sky130_fd_sc_hd__buf_1 _0631_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0123_),
    .X(_0124_)
);

sky130_fd_sc_hd__or2_4 _0632_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[31]),
    .B(_0124_),
    .X(_0125_)
);

sky130_fd_sc_hd__buf_1 _0633_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0105_),
    .X(_0126_)
);

sky130_fd_sc_hd__buf_1 _0634_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0126_),
    .X(_0127_)
);

sky130_fd_sc_hd__buf_1 _0635_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0127_),
    .X(_0128_)
);

sky130_fd_sc_hd__buf_1 _0636_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0111_),
    .X(_0129_)
);

sky130_fd_sc_hd__buf_1 _0637_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0129_),
    .X(_0130_)
);

sky130_fd_sc_hd__and2_4 _0638_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[31]),
    .B(_0130_),
    .X(_0131_)
);

sky130_fd_sc_hd__a21o_4 _0639_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[31]),
    .A2(_0128_),
    .B1(_0131_),
    .X(_0132_)
);

sky130_fd_sc_hd__and2_4 _0640_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[31]),
    .B(_0102_),
    .X(_0133_)
);

sky130_fd_sc_hd__a21o_4 _0641_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[31]),
    .A2(_0099_),
    .B1(_0133_),
    .X(_0134_)
);

sky130_fd_sc_hd__buf_1 _0642_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0093_),
    .X(_0135_)
);

sky130_fd_sc_hd__buf_1 _0643_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0108_),
    .X(_0136_)
);

sky130_fd_sc_hd__a21o_4 _0644_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[31]),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0137_)
);

sky130_fd_sc_hd__buf_1 _0645_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0116_),
    .X(_0138_)
);

sky130_fd_sc_hd__buf_1 _0646_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0087_),
    .X(_0139_)
);

sky130_fd_sc_hd__buf_1 _0647_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0139_),
    .X(_0140_)
);

sky130_fd_sc_hd__and2_4 _0648_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[31]),
    .B(_0140_),
    .X(_0141_)
);

sky130_fd_sc_hd__a21o_4 _0649_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[31]),
    .A2(_0138_),
    .B1(_0141_),
    .X(_0142_)
);

sky130_fd_sc_hd__or4_4 _0650_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0132_),
    .B(_0134_),
    .C(_0137_),
    .D(_0142_),
    .X(_0143_)
);

sky130_fd_sc_hd__and3_4 _0651_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .B(_0125_),
    .C(_0143_),
    .X(_0144_)
);

sky130_fd_sc_hd__nor3_4 _0652_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0120_),
    .C(_0144_),
    .Y(_0145_)
);

sky130_fd_sc_hd__or2_4 _0653_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[7]),
    .B(_0124_),
    .X(_0146_)
);

sky130_fd_sc_hd__and2_4 _0654_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[7]),
    .B(_0130_),
    .X(_0147_)
);

sky130_fd_sc_hd__a21o_4 _0655_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[7]),
    .A2(_0128_),
    .B1(_0147_),
    .X(_0148_)
);

sky130_fd_sc_hd__buf_1 _0656_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0098_),
    .X(_0149_)
);

sky130_fd_sc_hd__buf_1 _0657_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0149_),
    .X(_0150_)
);

sky130_fd_sc_hd__and2_4 _0658_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[7]),
    .B(_0102_),
    .X(_0151_)
);

sky130_fd_sc_hd__a21o_4 _0659_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[7]),
    .A2(_0150_),
    .B1(_0151_),
    .X(_0152_)
);

sky130_fd_sc_hd__a21o_4 _0660_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[7]),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0153_)
);

sky130_fd_sc_hd__buf_1 _0661_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0088_),
    .X(_0154_)
);

sky130_fd_sc_hd__buf_1 _0662_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0154_),
    .X(_0155_)
);

sky130_fd_sc_hd__and2_4 _0663_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[7]),
    .B(_0155_),
    .X(_0156_)
);

sky130_fd_sc_hd__a21o_4 _0664_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[7]),
    .A2(_0138_),
    .B1(_0156_),
    .X(_0157_)
);

sky130_fd_sc_hd__or4_4 _0665_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0148_),
    .B(_0152_),
    .C(_0153_),
    .D(_0157_),
    .X(_0158_)
);

sky130_fd_sc_hd__and3_4 _0666_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0077_),
    .B(_0146_),
    .C(_0158_),
    .X(_0159_)
);

sky130_fd_sc_hd__buf_1 _0667_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .X(_0160_)
);

sky130_fd_sc_hd__or2_4 _0668_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[23]),
    .B(_0124_),
    .X(_0161_)
);

sky130_fd_sc_hd__buf_1 _0669_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0111_),
    .X(_0162_)
);

sky130_fd_sc_hd__buf_1 _0670_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0162_),
    .X(_0163_)
);

sky130_fd_sc_hd__and2_4 _0671_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[23]),
    .B(_0163_),
    .X(_0164_)
);

sky130_fd_sc_hd__a21o_4 _0672_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[23]),
    .A2(_0128_),
    .B1(_0164_),
    .X(_0165_)
);

sky130_fd_sc_hd__and2_4 _0673_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[23]),
    .B(_0140_),
    .X(_0166_)
);

sky130_fd_sc_hd__a21o_4 _0674_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[23]),
    .A2(_0138_),
    .B1(_0166_),
    .X(_0167_)
);

sky130_fd_sc_hd__a21o_4 _0675_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[23]),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0168_)
);

sky130_fd_sc_hd__buf_1 _0676_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0098_),
    .X(_0169_)
);

sky130_fd_sc_hd__buf_1 _0677_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0169_),
    .X(_0170_)
);

sky130_fd_sc_hd__buf_1 _0678_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0101_),
    .X(_0171_)
);

sky130_fd_sc_hd__buf_1 _0679_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0171_),
    .X(_0172_)
);

sky130_fd_sc_hd__and2_4 _0680_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[23]),
    .B(_0172_),
    .X(_0173_)
);

sky130_fd_sc_hd__a21o_4 _0681_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[23]),
    .A2(_0170_),
    .B1(_0173_),
    .X(_0174_)
);

sky130_fd_sc_hd__or4_4 _0682_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0165_),
    .B(_0167_),
    .C(_0168_),
    .D(_0174_),
    .X(_0175_)
);

sky130_fd_sc_hd__and3_4 _0683_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .B(_0161_),
    .C(_0175_),
    .X(_0176_)
);

sky130_fd_sc_hd__nor3_4 _0684_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0069_),
    .B(_0159_),
    .C(_0176_),
    .Y(_0177_)
);

sky130_fd_sc_hd__nor3_4 _0685_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0064_),
    .B(_0145_),
    .C(_0177_),
    .Y(_0178_)
);

sky130_fd_sc_hd__or2_4 _0686_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[3]),
    .B(_0085_),
    .X(_0179_)
);

sky130_fd_sc_hd__and2_4 _0687_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[3]),
    .B(_0130_),
    .X(_0180_)
);

sky130_fd_sc_hd__a21o_4 _0688_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[3]),
    .A2(_0107_),
    .B1(_0180_),
    .X(_0181_)
);

sky130_fd_sc_hd__buf_1 _0689_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0116_),
    .X(_0182_)
);

sky130_fd_sc_hd__and2_4 _0690_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[3]),
    .B(_0140_),
    .X(_0183_)
);

sky130_fd_sc_hd__a21o_4 _0691_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[3]),
    .A2(_0182_),
    .B1(_0183_),
    .X(_0184_)
);

sky130_fd_sc_hd__buf_1 _0692_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0092_),
    .X(_0185_)
);

sky130_fd_sc_hd__a21o_4 _0693_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[3]),
    .A2(_0185_),
    .B1(_0109_),
    .X(_0186_)
);

sky130_fd_sc_hd__and2_4 _0694_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[3]),
    .B(_0172_),
    .X(_0187_)
);

sky130_fd_sc_hd__a21o_4 _0695_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[3]),
    .A2(_0150_),
    .B1(_0187_),
    .X(_0188_)
);

sky130_fd_sc_hd__or4_4 _0696_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0181_),
    .B(_0184_),
    .C(_0186_),
    .D(_0188_),
    .X(_0189_)
);

sky130_fd_sc_hd__and3_4 _0697_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0077_),
    .B(_0179_),
    .C(_0189_),
    .X(_0190_)
);

sky130_fd_sc_hd__or2_4 _0698_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[19]),
    .B(_0124_),
    .X(_0191_)
);

sky130_fd_sc_hd__and2_4 _0699_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[19]),
    .B(_0130_),
    .X(_0192_)
);

sky130_fd_sc_hd__a21o_4 _0700_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[19]),
    .A2(_0128_),
    .B1(_0192_),
    .X(_0193_)
);

sky130_fd_sc_hd__and2_4 _0701_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[19]),
    .B(_0172_),
    .X(_0194_)
);

sky130_fd_sc_hd__a21o_4 _0702_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[19]),
    .A2(_0150_),
    .B1(_0194_),
    .X(_0195_)
);

sky130_fd_sc_hd__a21o_4 _0703_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[19]),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0196_)
);

sky130_fd_sc_hd__buf_1 _0704_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0114_),
    .X(_0197_)
);

sky130_fd_sc_hd__buf_1 _0705_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0197_),
    .X(_0198_)
);

sky130_fd_sc_hd__buf_1 _0706_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0198_),
    .X(_0199_)
);

sky130_fd_sc_hd__and2_4 _0707_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[19]),
    .B(_0155_),
    .X(_0200_)
);

sky130_fd_sc_hd__a21o_4 _0708_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[19]),
    .A2(_0199_),
    .B1(_0200_),
    .X(_0201_)
);

sky130_fd_sc_hd__or4_4 _0709_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0193_),
    .B(_0195_),
    .C(_0196_),
    .D(_0201_),
    .X(_0202_)
);

sky130_fd_sc_hd__and3_4 _0710_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .B(_0191_),
    .C(_0202_),
    .X(_0203_)
);

sky130_fd_sc_hd__nor3_4 _0711_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0069_),
    .B(_0190_),
    .C(_0203_),
    .Y(_0204_)
);

sky130_fd_sc_hd__or2_4 _0712_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[27]),
    .B(_0124_),
    .X(_0205_)
);

sky130_fd_sc_hd__and2_4 _0713_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[27]),
    .B(_0163_),
    .X(_0206_)
);

sky130_fd_sc_hd__a21o_4 _0714_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[27]),
    .A2(_0128_),
    .B1(_0206_),
    .X(_0207_)
);

sky130_fd_sc_hd__and2_4 _0715_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[27]),
    .B(_0140_),
    .X(_0208_)
);

sky130_fd_sc_hd__a21o_4 _0716_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[27]),
    .A2(_0138_),
    .B1(_0208_),
    .X(_0209_)
);

sky130_fd_sc_hd__a21o_4 _0717_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[27]),
    .A2(_0135_),
    .B1(_0136_),
    .X(_0210_)
);

sky130_fd_sc_hd__and2_4 _0718_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[27]),
    .B(_0172_),
    .X(_0211_)
);

sky130_fd_sc_hd__a21o_4 _0719_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[27]),
    .A2(_0150_),
    .B1(_0211_),
    .X(_0212_)
);

sky130_fd_sc_hd__or4_4 _0720_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0207_),
    .B(_0209_),
    .C(_0210_),
    .D(_0212_),
    .X(_0213_)
);

sky130_fd_sc_hd__and3_4 _0721_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .B(_0205_),
    .C(_0213_),
    .X(_0214_)
);

sky130_fd_sc_hd__buf_1 _0722_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0085_),
    .X(_0215_)
);

sky130_fd_sc_hd__or2_4 _0723_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[11]),
    .B(_0215_),
    .X(_0216_)
);

sky130_fd_sc_hd__buf_1 _0724_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0106_),
    .X(_0217_)
);

sky130_fd_sc_hd__buf_1 _0725_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0217_),
    .X(_0218_)
);

sky130_fd_sc_hd__and2_4 _0726_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[11]),
    .B(_0163_),
    .X(_0219_)
);

sky130_fd_sc_hd__a21o_4 _0727_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[11]),
    .A2(_0218_),
    .B1(_0219_),
    .X(_0220_)
);

sky130_fd_sc_hd__and2_4 _0728_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[11]),
    .B(_0172_),
    .X(_0221_)
);

sky130_fd_sc_hd__a21o_4 _0729_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[11]),
    .A2(_0150_),
    .B1(_0221_),
    .X(_0222_)
);

sky130_fd_sc_hd__buf_1 _0730_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0092_),
    .X(_0223_)
);

sky130_fd_sc_hd__buf_1 _0731_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0223_),
    .X(_0224_)
);

sky130_fd_sc_hd__buf_1 _0732_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0108_),
    .X(_0225_)
);

sky130_fd_sc_hd__buf_1 _0733_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0225_),
    .X(_0226_)
);

sky130_fd_sc_hd__a21o_4 _0734_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[11]),
    .A2(_0224_),
    .B1(_0226_),
    .X(_0227_)
);

sky130_fd_sc_hd__and2_4 _0735_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[11]),
    .B(_0155_),
    .X(_0228_)
);

sky130_fd_sc_hd__a21o_4 _0736_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[11]),
    .A2(_0199_),
    .B1(_0228_),
    .X(_0229_)
);

sky130_fd_sc_hd__or4_4 _0737_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0220_),
    .B(_0222_),
    .C(_0227_),
    .D(_0229_),
    .X(_0230_)
);

sky130_fd_sc_hd__and3_4 _0738_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0017_),
    .B(_0216_),
    .C(_0230_),
    .X(_0231_)
);

sky130_fd_sc_hd__nor3_4 _0739_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0214_),
    .C(_0231_),
    .Y(_0232_)
);

sky130_fd_sc_hd__nor3_4 _0740_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[2]),
    .B(_0204_),
    .C(_0232_),
    .Y(_0233_)
);

sky130_fd_sc_hd__or2_4 _0741_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[5]),
    .B(_0215_),
    .X(_0234_)
);

sky130_fd_sc_hd__and2_4 _0742_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[5]),
    .B(_0163_),
    .X(_0235_)
);

sky130_fd_sc_hd__a21o_4 _0743_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[5]),
    .A2(_0218_),
    .B1(_0235_),
    .X(_0236_)
);

sky130_fd_sc_hd__and2_4 _0744_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[5]),
    .B(_0155_),
    .X(_0237_)
);

sky130_fd_sc_hd__a21o_4 _0745_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[5]),
    .A2(_0138_),
    .B1(_0237_),
    .X(_0238_)
);

sky130_fd_sc_hd__a21o_4 _0746_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[5]),
    .A2(_0224_),
    .B1(_0226_),
    .X(_0239_)
);

sky130_fd_sc_hd__buf_1 _0747_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0101_),
    .X(_0240_)
);

sky130_fd_sc_hd__buf_1 _0748_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0240_),
    .X(_0241_)
);

sky130_fd_sc_hd__and2_4 _0749_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[5]),
    .B(_0241_),
    .X(_0242_)
);

sky130_fd_sc_hd__a21o_4 _0750_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[5]),
    .A2(_0170_),
    .B1(_0242_),
    .X(_0243_)
);

sky130_fd_sc_hd__or4_4 _0751_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0236_),
    .B(_0238_),
    .C(_0239_),
    .D(_0243_),
    .X(_0244_)
);

sky130_fd_sc_hd__and3_4 _0752_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0017_),
    .B(_0234_),
    .C(_0244_),
    .X(_0245_)
);

sky130_fd_sc_hd__or2_4 _0753_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[21]),
    .B(_0215_),
    .X(_0246_)
);

sky130_fd_sc_hd__and2_4 _0754_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[21]),
    .B(_0163_),
    .X(_0247_)
);

sky130_fd_sc_hd__a21o_4 _0755_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[21]),
    .A2(_0218_),
    .B1(_0247_),
    .X(_0248_)
);

sky130_fd_sc_hd__and2_4 _0756_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[21]),
    .B(_0241_),
    .X(_0249_)
);

sky130_fd_sc_hd__a21o_4 _0757_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[21]),
    .A2(_0170_),
    .B1(_0249_),
    .X(_0250_)
);

sky130_fd_sc_hd__a21o_4 _0758_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[21]),
    .A2(_0224_),
    .B1(_0226_),
    .X(_0251_)
);

sky130_fd_sc_hd__and2_4 _0759_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[21]),
    .B(_0090_),
    .X(_0252_)
);

sky130_fd_sc_hd__a21o_4 _0760_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[21]),
    .A2(_0199_),
    .B1(_0252_),
    .X(_0253_)
);

sky130_fd_sc_hd__or4_4 _0761_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0248_),
    .B(_0250_),
    .C(_0251_),
    .D(_0253_),
    .X(_0254_)
);

sky130_fd_sc_hd__and3_4 _0762_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .B(_0246_),
    .C(_0254_),
    .X(_0255_)
);

sky130_fd_sc_hd__nor3_4 _0763_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0069_),
    .B(_0245_),
    .C(_0255_),
    .Y(_0256_)
);

sky130_fd_sc_hd__or2_4 _0764_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[29]),
    .B(_0215_),
    .X(_0257_)
);

sky130_fd_sc_hd__and2_4 _0765_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[29]),
    .B(_0113_),
    .X(_0258_)
);

sky130_fd_sc_hd__a21o_4 _0766_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[29]),
    .A2(_0218_),
    .B1(_0258_),
    .X(_0259_)
);

sky130_fd_sc_hd__and2_4 _0767_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[29]),
    .B(_0241_),
    .X(_0260_)
);

sky130_fd_sc_hd__a21o_4 _0768_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[29]),
    .A2(_0170_),
    .B1(_0260_),
    .X(_0261_)
);

sky130_fd_sc_hd__a21o_4 _0769_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[29]),
    .A2(_0224_),
    .B1(_0226_),
    .X(_0262_)
);

sky130_fd_sc_hd__and2_4 _0770_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[29]),
    .B(_0090_),
    .X(_0263_)
);

sky130_fd_sc_hd__a21o_4 _0771_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[29]),
    .A2(_0199_),
    .B1(_0263_),
    .X(_0264_)
);

sky130_fd_sc_hd__or4_4 _0772_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0259_),
    .B(_0261_),
    .C(_0262_),
    .D(_0264_),
    .X(_0265_)
);

sky130_fd_sc_hd__and3_4 _0773_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0160_),
    .B(_0257_),
    .C(_0265_),
    .X(_0266_)
);

sky130_fd_sc_hd__or2_4 _0774_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[13]),
    .B(_0215_),
    .X(_0267_)
);

sky130_fd_sc_hd__and2_4 _0775_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[13]),
    .B(_0113_),
    .X(_0268_)
);

sky130_fd_sc_hd__a21o_4 _0776_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[13]),
    .A2(_0218_),
    .B1(_0268_),
    .X(_0269_)
);

sky130_fd_sc_hd__and2_4 _0777_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[13]),
    .B(_0090_),
    .X(_0270_)
);

sky130_fd_sc_hd__a21o_4 _0778_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[13]),
    .A2(_0199_),
    .B1(_0270_),
    .X(_0271_)
);

sky130_fd_sc_hd__a21o_4 _0779_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[13]),
    .A2(_0224_),
    .B1(_0226_),
    .X(_0272_)
);

sky130_fd_sc_hd__and2_4 _0780_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[13]),
    .B(_0241_),
    .X(_0273_)
);

sky130_fd_sc_hd__a21o_4 _0781_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[13]),
    .A2(_0170_),
    .B1(_0273_),
    .X(_0274_)
);

sky130_fd_sc_hd__or4_4 _0782_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0269_),
    .B(_0271_),
    .C(_0272_),
    .D(_0274_),
    .X(_0275_)
);

sky130_fd_sc_hd__and3_4 _0783_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0017_),
    .B(_0267_),
    .C(_0275_),
    .X(_0276_)
);

sky130_fd_sc_hd__nor3_4 _0784_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0266_),
    .C(_0276_),
    .Y(_0277_)
);

sky130_fd_sc_hd__nor3_4 _0785_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0064_),
    .B(_0256_),
    .C(_0277_),
    .Y(_0278_)
);

sky130_fd_sc_hd__or2_4 _0786_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[9]),
    .B(_0123_),
    .X(_0279_)
);

sky130_fd_sc_hd__and2_4 _0787_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[9]),
    .B(_0092_),
    .X(_0280_)
);

sky130_fd_sc_hd__a21o_4 _0788_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[9]),
    .A2(_0155_),
    .B1(_0280_),
    .X(_0281_)
);

sky130_fd_sc_hd__buf_1 _0789_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0100_),
    .X(_0282_)
);

sky130_fd_sc_hd__and2_4 _0790_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[9]),
    .B(_0282_),
    .X(_0283_)
);

sky130_fd_sc_hd__a21o_4 _0791_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[9]),
    .A2(_0149_),
    .B1(_0283_),
    .X(_0284_)
);

sky130_fd_sc_hd__buf_1 _0792_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0108_),
    .X(_0285_)
);

sky130_fd_sc_hd__a21o_4 _0793_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[9]),
    .A2(_0217_),
    .B1(_0285_),
    .X(_0286_)
);

sky130_fd_sc_hd__and2_4 _0794_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[9]),
    .B(_0197_),
    .X(_0287_)
);

sky130_fd_sc_hd__a21o_4 _0795_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[9]),
    .A2(_0113_),
    .B1(_0287_),
    .X(_0288_)
);

sky130_fd_sc_hd__or4_4 _0796_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0281_),
    .B(_0284_),
    .C(_0286_),
    .D(_0288_),
    .X(_0289_)
);

sky130_fd_sc_hd__and3_4 _0797_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0016_),
    .B(_0279_),
    .C(_0289_),
    .X(_0290_)
);

sky130_fd_sc_hd__buf_1 _0798_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0084_),
    .X(_0291_)
);

sky130_fd_sc_hd__or2_4 _0799_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[25]),
    .B(_0291_),
    .X(_0292_)
);

sky130_fd_sc_hd__buf_1 _0800_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0111_),
    .X(_0293_)
);

sky130_fd_sc_hd__and2_4 _0801_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[25]),
    .B(_0293_),
    .X(_0294_)
);

sky130_fd_sc_hd__a21o_4 _0802_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[25]),
    .A2(_0217_),
    .B1(_0294_),
    .X(_0295_)
);

sky130_fd_sc_hd__and2_4 _0803_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[25]),
    .B(_0240_),
    .X(_0296_)
);

sky130_fd_sc_hd__a21o_4 _0804_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[25]),
    .A2(_0169_),
    .B1(_0296_),
    .X(_0297_)
);

sky130_fd_sc_hd__a21o_4 _0805_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[25]),
    .A2(_0223_),
    .B1(_0225_),
    .X(_0298_)
);

sky130_fd_sc_hd__and2_4 _0806_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[25]),
    .B(_0089_),
    .X(_0299_)
);

sky130_fd_sc_hd__a21o_4 _0807_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[25]),
    .A2(_0182_),
    .B1(_0299_),
    .X(_0300_)
);

sky130_fd_sc_hd__or4_4 _0808_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0295_),
    .B(_0297_),
    .C(_0298_),
    .D(_0300_),
    .X(_0301_)
);

sky130_fd_sc_hd__and3_4 _0809_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .B(_0292_),
    .C(_0301_),
    .X(_0302_)
);

sky130_fd_sc_hd__nor3_4 _0810_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0019_),
    .B(_0290_),
    .C(_0302_),
    .Y(_0303_)
);

sky130_fd_sc_hd__or2_4 _0811_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[1]),
    .B(_0291_),
    .X(_0304_)
);

sky130_fd_sc_hd__and2_4 _0812_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[1]),
    .B(_0293_),
    .X(_0305_)
);

sky130_fd_sc_hd__a21o_4 _0813_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[1]),
    .A2(_0107_),
    .B1(_0305_),
    .X(_0306_)
);

sky130_fd_sc_hd__and2_4 _0814_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[1]),
    .B(_0154_),
    .X(_0307_)
);

sky130_fd_sc_hd__a21o_4 _0815_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[1]),
    .A2(_0198_),
    .B1(_0307_),
    .X(_0308_)
);

sky130_fd_sc_hd__a21o_4 _0816_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[1]),
    .A2(_0185_),
    .B1(_0109_),
    .X(_0309_)
);

sky130_fd_sc_hd__and2_4 _0817_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[1]),
    .B(_0102_),
    .X(_0310_)
);

sky130_fd_sc_hd__a21o_4 _0818_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[1]),
    .A2(_0099_),
    .B1(_0310_),
    .X(_0311_)
);

sky130_fd_sc_hd__or4_4 _0819_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0306_),
    .B(_0308_),
    .C(_0309_),
    .D(_0311_),
    .X(_0312_)
);

sky130_fd_sc_hd__and3_4 _0820_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0077_),
    .B(_0304_),
    .C(_0312_),
    .X(_0313_)
);

sky130_fd_sc_hd__or2_4 _0821_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[17]),
    .B(_0085_),
    .X(_0314_)
);

sky130_fd_sc_hd__and2_4 _0822_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[17]),
    .B(_0293_),
    .X(_0315_)
);

sky130_fd_sc_hd__a21o_4 _0823_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[17]),
    .A2(_0107_),
    .B1(_0315_),
    .X(_0316_)
);

sky130_fd_sc_hd__and2_4 _0824_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[17]),
    .B(_0102_),
    .X(_0317_)
);

sky130_fd_sc_hd__a21o_4 _0825_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[17]),
    .A2(_0099_),
    .B1(_0317_),
    .X(_0318_)
);

sky130_fd_sc_hd__a21o_4 _0826_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[17]),
    .A2(_0185_),
    .B1(_0109_),
    .X(_0319_)
);

sky130_fd_sc_hd__and2_4 _0827_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[17]),
    .B(_0140_),
    .X(_0320_)
);

sky130_fd_sc_hd__a21o_4 _0828_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[17]),
    .A2(_0182_),
    .B1(_0320_),
    .X(_0321_)
);

sky130_fd_sc_hd__or4_4 _0829_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0316_),
    .B(_0318_),
    .C(_0319_),
    .D(_0321_),
    .X(_0322_)
);

sky130_fd_sc_hd__and3_4 _0830_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .B(_0314_),
    .C(_0322_),
    .X(_0323_)
);

sky130_fd_sc_hd__nor3_4 _0831_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0069_),
    .B(_0313_),
    .C(_0323_),
    .Y(_0324_)
);

sky130_fd_sc_hd__nor3_4 _0832_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[2]),
    .B(_0303_),
    .C(_0324_),
    .Y(_0325_)
);

sky130_fd_sc_hd__or2_4 _0833_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[1]),
    .B(_0325_),
    .X(_0326_)
);

sky130_fd_sc_hd__o32ai_4 _0834_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0022_),
    .A2(_0178_),
    .A3(_0233_),
    .B1(_0278_),
    .B2(_0326_),
    .Y(_0327_)
);

sky130_fd_sc_hd__and2_4 _0835_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[0]),
    .B(_0327_),
    .X(_0328_)
);

sky130_fd_sc_hd__or2_4 _0836_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[10]),
    .B(_0083_),
    .X(_0329_)
);

sky130_fd_sc_hd__and2_4 _0837_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[10]),
    .B(_0091_),
    .X(_0330_)
);

sky130_fd_sc_hd__a21o_4 _0838_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[10]),
    .A2(_0129_),
    .B1(_0330_),
    .X(_0331_)
);

sky130_fd_sc_hd__and2_4 _0839_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[10]),
    .B(_0087_),
    .X(_0332_)
);

sky130_fd_sc_hd__a21o_4 _0840_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[10]),
    .A2(_0115_),
    .B1(_0332_),
    .X(_0333_)
);

sky130_fd_sc_hd__a21o_4 _0841_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[10]),
    .A2(_0097_),
    .B1(_0081_),
    .X(_0334_)
);

sky130_fd_sc_hd__and2_4 _0842_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN3[10]),
    .B(_0105_),
    .X(_0335_)
);

sky130_fd_sc_hd__a21o_4 _0843_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[10]),
    .A2(_0282_),
    .B1(_0335_),
    .X(_0336_)
);

sky130_fd_sc_hd__or4_4 _0844_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0331_),
    .B(_0333_),
    .C(_0334_),
    .D(_0336_),
    .X(_0337_)
);

sky130_fd_sc_hd__and3_4 _0845_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0015_),
    .B(_0329_),
    .C(_0337_),
    .X(_0338_)
);

sky130_fd_sc_hd__or2_4 _0846_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[26]),
    .B(_0083_),
    .X(_0339_)
);

sky130_fd_sc_hd__and2_4 _0847_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[26]),
    .B(_0091_),
    .X(_0340_)
);

sky130_fd_sc_hd__a21o_4 _0848_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[26]),
    .A2(_0101_),
    .B1(_0340_),
    .X(_0341_)
);

sky130_fd_sc_hd__and2_4 _0849_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[26]),
    .B(_0087_),
    .X(_0342_)
);

sky130_fd_sc_hd__a21o_4 _0850_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[26]),
    .A2(_0115_),
    .B1(_0342_),
    .X(_0343_)
);

sky130_fd_sc_hd__a21o_4 _0851_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[26]),
    .A2(_0105_),
    .B1(_0081_),
    .X(_0344_)
);

sky130_fd_sc_hd__and2_4 _0852_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN8[26]),
    .B(_0096_),
    .X(_0345_)
);

sky130_fd_sc_hd__a21o_4 _0853_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[26]),
    .A2(_0129_),
    .B1(_0345_),
    .X(_0346_)
);

sky130_fd_sc_hd__or4_4 _0854_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0341_),
    .B(_0343_),
    .C(_0344_),
    .D(_0346_),
    .X(_0347_)
);

sky130_fd_sc_hd__and3_4 _0855_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[4]),
    .B(_0339_),
    .C(_0347_),
    .X(_0348_)
);

sky130_fd_sc_hd__or3_4 _0856_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0018_),
    .B(_0338_),
    .C(_0348_),
    .X(_0349_)
);

sky130_fd_sc_hd__buf_1 _0857_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0083_),
    .X(_0350_)
);

sky130_fd_sc_hd__or2_4 _0858_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[18]),
    .B(_0350_),
    .X(_0351_)
);

sky130_fd_sc_hd__buf_1 _0859_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0091_),
    .X(_0352_)
);

sky130_fd_sc_hd__and2_4 _0860_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[18]),
    .B(_0352_),
    .X(_0353_)
);

sky130_fd_sc_hd__a21o_4 _0861_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[18]),
    .A2(_0282_),
    .B1(_0353_),
    .X(_0354_)
);

sky130_fd_sc_hd__and2_4 _0862_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[18]),
    .B(_0088_),
    .X(_0355_)
);

sky130_fd_sc_hd__a21o_4 _0863_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[18]),
    .A2(_0115_),
    .B1(_0355_),
    .X(_0356_)
);

sky130_fd_sc_hd__a21o_4 _0864_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[18]),
    .A2(_0126_),
    .B1(_0081_),
    .X(_0357_)
);

sky130_fd_sc_hd__and2_4 _0865_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN8[18]),
    .B(_0096_),
    .X(_0358_)
);

sky130_fd_sc_hd__a21o_4 _0866_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[18]),
    .A2(_0129_),
    .B1(_0358_),
    .X(_0359_)
);

sky130_fd_sc_hd__or4_4 _0867_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0354_),
    .B(_0356_),
    .C(_0357_),
    .D(_0359_),
    .X(_0360_)
);

sky130_fd_sc_hd__and3_4 _0868_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[4]),
    .B(_0351_),
    .C(_0360_),
    .X(_0361_)
);

sky130_fd_sc_hd__or2_4 _0869_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[2]),
    .B(_0350_),
    .X(_0362_)
);

sky130_fd_sc_hd__and2_4 _0870_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[2]),
    .B(_0352_),
    .X(_0363_)
);

sky130_fd_sc_hd__a21o_4 _0871_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[2]),
    .A2(_0139_),
    .B1(_0363_),
    .X(_0364_)
);

sky130_fd_sc_hd__and2_4 _0872_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[2]),
    .B(_0100_),
    .X(_0365_)
);

sky130_fd_sc_hd__a21o_4 _0873_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[2]),
    .A2(_0097_),
    .B1(_0365_),
    .X(_0366_)
);

sky130_fd_sc_hd__a21o_4 _0874_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[2]),
    .A2(_0126_),
    .B1(_0082_),
    .X(_0367_)
);

sky130_fd_sc_hd__and2_4 _0875_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[2]),
    .B(_0114_),
    .X(_0368_)
);

sky130_fd_sc_hd__a21o_4 _0876_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[2]),
    .A2(_0129_),
    .B1(_0368_),
    .X(_0369_)
);

sky130_fd_sc_hd__or4_4 _0877_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0364_),
    .B(_0366_),
    .C(_0367_),
    .D(_0369_),
    .X(_0370_)
);

sky130_fd_sc_hd__and3_4 _0878_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0015_),
    .B(_0362_),
    .C(_0370_),
    .X(_0371_)
);

sky130_fd_sc_hd__or3_4 _0879_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0068_),
    .B(_0361_),
    .C(_0371_),
    .X(_0372_)
);

sky130_fd_sc_hd__or2_4 _0880_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[30]),
    .B(_0350_),
    .X(_0373_)
);

sky130_fd_sc_hd__and2_4 _0881_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[30]),
    .B(_0352_),
    .X(_0374_)
);

sky130_fd_sc_hd__a21o_4 _0882_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[30]),
    .A2(_0282_),
    .B1(_0374_),
    .X(_0375_)
);

sky130_fd_sc_hd__and2_4 _0883_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[30]),
    .B(_0088_),
    .X(_0376_)
);

sky130_fd_sc_hd__a21o_4 _0884_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[30]),
    .A2(_0197_),
    .B1(_0376_),
    .X(_0377_)
);

sky130_fd_sc_hd__a21o_4 _0885_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[30]),
    .A2(_0126_),
    .B1(_0082_),
    .X(_0378_)
);

sky130_fd_sc_hd__and2_4 _0886_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN8[30]),
    .B(_0096_),
    .X(_0379_)
);

sky130_fd_sc_hd__a21o_4 _0887_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[30]),
    .A2(_0112_),
    .B1(_0379_),
    .X(_0380_)
);

sky130_fd_sc_hd__or4_4 _0888_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0375_),
    .B(_0377_),
    .C(_0378_),
    .D(_0380_),
    .X(_0381_)
);

sky130_fd_sc_hd__and3_4 _0889_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[4]),
    .B(_0373_),
    .C(_0381_),
    .X(_0382_)
);

sky130_fd_sc_hd__or2_4 _0890_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[14]),
    .B(_0350_),
    .X(_0383_)
);

sky130_fd_sc_hd__and2_4 _0891_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[14]),
    .B(_0352_),
    .X(_0384_)
);

sky130_fd_sc_hd__a21o_4 _0892_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[14]),
    .A2(_0139_),
    .B1(_0384_),
    .X(_0385_)
);

sky130_fd_sc_hd__and2_4 _0893_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[14]),
    .B(_0100_),
    .X(_0386_)
);

sky130_fd_sc_hd__a21o_4 _0894_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[14]),
    .A2(_0097_),
    .B1(_0386_),
    .X(_0387_)
);

sky130_fd_sc_hd__a21o_4 _0895_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[14]),
    .A2(_0126_),
    .B1(_0082_),
    .X(_0388_)
);

sky130_fd_sc_hd__and2_4 _0896_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[14]),
    .B(_0114_),
    .X(_0389_)
);

sky130_fd_sc_hd__a21o_4 _0897_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[14]),
    .A2(_0112_),
    .B1(_0389_),
    .X(_0390_)
);

sky130_fd_sc_hd__or4_4 _0898_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0385_),
    .B(_0387_),
    .C(_0388_),
    .D(_0390_),
    .X(_0391_)
);

sky130_fd_sc_hd__and3_4 _0899_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0015_),
    .B(_0383_),
    .C(_0391_),
    .X(_0392_)
);

sky130_fd_sc_hd__or3_4 _0900_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0019_),
    .B(_0382_),
    .C(_0392_),
    .X(_0393_)
);

sky130_fd_sc_hd__or2_4 _0901_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[22]),
    .B(_0350_),
    .X(_0394_)
);

sky130_fd_sc_hd__and2_4 _0902_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[22]),
    .B(_0352_),
    .X(_0395_)
);

sky130_fd_sc_hd__a21o_4 _0903_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[22]),
    .A2(_0282_),
    .B1(_0395_),
    .X(_0396_)
);

sky130_fd_sc_hd__and2_4 _0904_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[22]),
    .B(_0088_),
    .X(_0397_)
);

sky130_fd_sc_hd__a21o_4 _0905_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[22]),
    .A2(_0197_),
    .B1(_0397_),
    .X(_0398_)
);

sky130_fd_sc_hd__a21o_4 _0906_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[22]),
    .A2(_0106_),
    .B1(_0082_),
    .X(_0399_)
);

sky130_fd_sc_hd__and2_4 _0907_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN8[22]),
    .B(_0097_),
    .X(_0400_)
);

sky130_fd_sc_hd__a21o_4 _0908_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[22]),
    .A2(_0293_),
    .B1(_0400_),
    .X(_0401_)
);

sky130_fd_sc_hd__or4_4 _0909_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0396_),
    .B(_0398_),
    .C(_0399_),
    .D(_0401_),
    .X(_0402_)
);

sky130_fd_sc_hd__and3_4 _0910_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0121_),
    .B(_0394_),
    .C(_0402_),
    .X(_0403_)
);

sky130_fd_sc_hd__and2_4 _0911_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN4[6]),
    .B(_0092_),
    .X(_0404_)
);

sky130_fd_sc_hd__a21o_4 _0912_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[6]),
    .A2(_0154_),
    .B1(_0404_),
    .X(_0405_)
);

sky130_fd_sc_hd__and2_4 _0913_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[6]),
    .B(_0101_),
    .X(_0406_)
);

sky130_fd_sc_hd__a21o_4 _0914_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[6]),
    .A2(_0098_),
    .B1(_0406_),
    .X(_0407_)
);

sky130_fd_sc_hd__a21o_4 _0915_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[6]),
    .A2(_0106_),
    .B1(_0108_),
    .X(_0408_)
);

sky130_fd_sc_hd__and2_4 _0916_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[6]),
    .B(_0115_),
    .X(_0409_)
);

sky130_fd_sc_hd__a21o_4 _0917_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[6]),
    .A2(_0130_),
    .B1(_0409_),
    .X(_0410_)
);

sky130_fd_sc_hd__or4_4 _0918_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0405_),
    .B(_0407_),
    .C(_0408_),
    .D(_0410_),
    .X(_0411_)
);

sky130_fd_sc_hd__o21a_4 _0919_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN1[6]),
    .A2(_0084_),
    .B1(_0014_),
    .X(_0412_)
);

sky130_fd_sc_hd__a21o_4 _0920_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0411_),
    .A2(_0412_),
    .B1(_0068_),
    .X(_0413_)
);

sky130_fd_sc_hd__o21a_4 _0921_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0403_),
    .A2(_0413_),
    .B1(COUNT[2]),
    .X(_0414_)
);

sky130_fd_sc_hd__a32o_4 _0922_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0020_),
    .A2(_0349_),
    .A3(_0372_),
    .B1(_0393_),
    .B2(_0414_),
    .X(_0415_)
);

sky130_fd_sc_hd__and2_4 _0923_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[1]),
    .B(_0415_),
    .X(_0416_)
);

sky130_fd_sc_hd__or2_4 _0924_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[0]),
    .B(_0084_),
    .X(_0417_)
);

sky130_fd_sc_hd__and2_4 _0925_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[0]),
    .B(_0112_),
    .X(_0418_)
);

sky130_fd_sc_hd__a21o_4 _0926_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[0]),
    .A2(_0127_),
    .B1(_0418_),
    .X(_0419_)
);

sky130_fd_sc_hd__and2_4 _0927_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[0]),
    .B(_0139_),
    .X(_0420_)
);

sky130_fd_sc_hd__a21o_4 _0928_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[0]),
    .A2(_0116_),
    .B1(_0420_),
    .X(_0421_)
);

sky130_fd_sc_hd__a21o_4 _0929_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[0]),
    .A2(_0093_),
    .B1(_0285_),
    .X(_0422_)
);

sky130_fd_sc_hd__and2_4 _0930_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[0]),
    .B(_0171_),
    .X(_0423_)
);

sky130_fd_sc_hd__a21o_4 _0931_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[0]),
    .A2(_0149_),
    .B1(_0423_),
    .X(_0424_)
);

sky130_fd_sc_hd__or4_4 _0932_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0419_),
    .B(_0421_),
    .C(_0422_),
    .D(_0424_),
    .X(_0425_)
);

sky130_fd_sc_hd__and3_4 _0933_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0016_),
    .B(_0417_),
    .C(_0425_),
    .X(_0426_)
);

sky130_fd_sc_hd__or2_4 _0934_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[16]),
    .B(_0123_),
    .X(_0427_)
);

sky130_fd_sc_hd__and2_4 _0935_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[16]),
    .B(_0162_),
    .X(_0428_)
);

sky130_fd_sc_hd__a21o_4 _0936_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[16]),
    .A2(_0127_),
    .B1(_0428_),
    .X(_0429_)
);

sky130_fd_sc_hd__and2_4 _0937_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[16]),
    .B(_0171_),
    .X(_0430_)
);

sky130_fd_sc_hd__a21o_4 _0938_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[16]),
    .A2(_0149_),
    .B1(_0430_),
    .X(_0431_)
);

sky130_fd_sc_hd__a21o_4 _0939_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[16]),
    .A2(_0093_),
    .B1(_0285_),
    .X(_0432_)
);

sky130_fd_sc_hd__and2_4 _0940_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[16]),
    .B(_0154_),
    .X(_0433_)
);

sky130_fd_sc_hd__a21o_4 _0941_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[16]),
    .A2(_0198_),
    .B1(_0433_),
    .X(_0434_)
);

sky130_fd_sc_hd__or4_4 _0942_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0429_),
    .B(_0431_),
    .C(_0432_),
    .D(_0434_),
    .X(_0435_)
);

sky130_fd_sc_hd__and3_4 _0943_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0121_),
    .B(_0427_),
    .C(_0435_),
    .X(_0436_)
);

sky130_fd_sc_hd__nor3_4 _0944_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0068_),
    .B(_0426_),
    .C(_0436_),
    .Y(_0437_)
);

sky130_fd_sc_hd__or2_4 _0945_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[24]),
    .B(_0123_),
    .X(_0438_)
);

sky130_fd_sc_hd__and2_4 _0946_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[24]),
    .B(_0162_),
    .X(_0439_)
);

sky130_fd_sc_hd__a21o_4 _0947_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[24]),
    .A2(_0127_),
    .B1(_0439_),
    .X(_0440_)
);

sky130_fd_sc_hd__and2_4 _0948_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[24]),
    .B(_0154_),
    .X(_0441_)
);

sky130_fd_sc_hd__a21o_4 _0949_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[24]),
    .A2(_0198_),
    .B1(_0441_),
    .X(_0442_)
);

sky130_fd_sc_hd__a21o_4 _0950_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[24]),
    .A2(_0223_),
    .B1(_0285_),
    .X(_0443_)
);

sky130_fd_sc_hd__and2_4 _0951_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[24]),
    .B(_0240_),
    .X(_0444_)
);

sky130_fd_sc_hd__a21o_4 _0952_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[24]),
    .A2(_0099_),
    .B1(_0444_),
    .X(_0445_)
);

sky130_fd_sc_hd__or4_4 _0953_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0440_),
    .B(_0442_),
    .C(_0443_),
    .D(_0445_),
    .X(_0446_)
);

sky130_fd_sc_hd__and3_4 _0954_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0121_),
    .B(_0438_),
    .C(_0446_),
    .X(_0447_)
);

sky130_fd_sc_hd__or2_4 _0955_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[8]),
    .B(_0291_),
    .X(_0448_)
);

sky130_fd_sc_hd__and2_4 _0956_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[8]),
    .B(_0293_),
    .X(_0449_)
);

sky130_fd_sc_hd__a21o_4 _0957_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[8]),
    .A2(_0107_),
    .B1(_0449_),
    .X(_0450_)
);

sky130_fd_sc_hd__and2_4 _0958_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[8]),
    .B(_0240_),
    .X(_0451_)
);

sky130_fd_sc_hd__a21o_4 _0959_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[8]),
    .A2(_0169_),
    .B1(_0451_),
    .X(_0452_)
);

sky130_fd_sc_hd__a21o_4 _0960_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[8]),
    .A2(_0185_),
    .B1(_0225_),
    .X(_0453_)
);

sky130_fd_sc_hd__and2_4 _0961_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[8]),
    .B(_0089_),
    .X(_0454_)
);

sky130_fd_sc_hd__a21o_4 _0962_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[8]),
    .A2(_0182_),
    .B1(_0454_),
    .X(_0455_)
);

sky130_fd_sc_hd__or4_4 _0963_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0450_),
    .B(_0452_),
    .C(_0453_),
    .D(_0455_),
    .X(_0456_)
);

sky130_fd_sc_hd__and3_4 _0964_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0077_),
    .B(_0448_),
    .C(_0456_),
    .X(_0457_)
);

sky130_fd_sc_hd__nor3_4 _0965_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0072_),
    .B(_0447_),
    .C(_0457_),
    .Y(_0458_)
);

sky130_fd_sc_hd__nor3_4 _0966_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[2]),
    .B(_0437_),
    .C(_0458_),
    .Y(_0459_)
);

sky130_fd_sc_hd__or2_4 _0967_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[28]),
    .B(_0123_),
    .X(_0460_)
);

sky130_fd_sc_hd__and2_4 _0968_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[28]),
    .B(_0112_),
    .X(_0461_)
);

sky130_fd_sc_hd__a21o_4 _0969_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[28]),
    .A2(_0127_),
    .B1(_0461_),
    .X(_0462_)
);

sky130_fd_sc_hd__and2_4 _0970_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[28]),
    .B(_0139_),
    .X(_0463_)
);

sky130_fd_sc_hd__a21o_4 _0971_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[28]),
    .A2(_0116_),
    .B1(_0463_),
    .X(_0464_)
);

sky130_fd_sc_hd__a21o_4 _0972_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[28]),
    .A2(_0093_),
    .B1(_0285_),
    .X(_0465_)
);

sky130_fd_sc_hd__and2_4 _0973_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[28]),
    .B(_0240_),
    .X(_0466_)
);

sky130_fd_sc_hd__a21o_4 _0974_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[28]),
    .A2(_0169_),
    .B1(_0466_),
    .X(_0467_)
);

sky130_fd_sc_hd__or4_4 _0975_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0462_),
    .B(_0464_),
    .C(_0465_),
    .D(_0467_),
    .X(_0468_)
);

sky130_fd_sc_hd__and3_4 _0976_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0121_),
    .B(_0460_),
    .C(_0468_),
    .X(_0469_)
);

sky130_fd_sc_hd__or2_4 _0977_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[12]),
    .B(_0291_),
    .X(_0470_)
);

sky130_fd_sc_hd__and2_4 _0978_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[12]),
    .B(_0162_),
    .X(_0471_)
);

sky130_fd_sc_hd__a21o_4 _0979_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[12]),
    .A2(_0217_),
    .B1(_0471_),
    .X(_0472_)
);

sky130_fd_sc_hd__and2_4 _0980_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[12]),
    .B(_0171_),
    .X(_0473_)
);

sky130_fd_sc_hd__a21o_4 _0981_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[12]),
    .A2(_0149_),
    .B1(_0473_),
    .X(_0474_)
);

sky130_fd_sc_hd__a21o_4 _0982_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[12]),
    .A2(_0223_),
    .B1(_0225_),
    .X(_0475_)
);

sky130_fd_sc_hd__and2_4 _0983_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[12]),
    .B(_0089_),
    .X(_0476_)
);

sky130_fd_sc_hd__a21o_4 _0984_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[12]),
    .A2(_0198_),
    .B1(_0476_),
    .X(_0477_)
);

sky130_fd_sc_hd__or4_4 _0985_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0472_),
    .B(_0474_),
    .C(_0475_),
    .D(_0477_),
    .X(_0478_)
);

sky130_fd_sc_hd__and3_4 _0986_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0016_),
    .B(_0470_),
    .C(_0478_),
    .X(_0479_)
);

sky130_fd_sc_hd__nor3_4 _0987_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0019_),
    .B(_0469_),
    .C(_0479_),
    .Y(_0480_)
);

sky130_fd_sc_hd__or2_4 _0988_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[4]),
    .B(_0291_),
    .X(_0481_)
);

sky130_fd_sc_hd__and2_4 _0989_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN2[4]),
    .B(_0162_),
    .X(_0482_)
);

sky130_fd_sc_hd__a21o_4 _0990_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN3[4]),
    .A2(_0217_),
    .B1(_0482_),
    .X(_0483_)
);

sky130_fd_sc_hd__and2_4 _0991_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN5[4]),
    .B(_0171_),
    .X(_0484_)
);

sky130_fd_sc_hd__a21o_4 _0992_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN8[4]),
    .A2(_0169_),
    .B1(_0484_),
    .X(_0485_)
);

sky130_fd_sc_hd__a21o_4 _0993_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[4]),
    .A2(_0223_),
    .B1(_0225_),
    .X(_0486_)
);

sky130_fd_sc_hd__and2_4 _0994_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN6[4]),
    .B(_0089_),
    .X(_0487_)
);

sky130_fd_sc_hd__a21o_4 _0995_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN7[4]),
    .A2(_0182_),
    .B1(_0487_),
    .X(_0488_)
);

sky130_fd_sc_hd__or4_4 _0996_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0483_),
    .B(_0485_),
    .C(_0486_),
    .D(_0488_),
    .X(_0489_)
);

sky130_fd_sc_hd__and3_4 _0997_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0016_),
    .B(_0481_),
    .C(_0489_),
    .X(_0490_)
);

sky130_fd_sc_hd__or2_4 _0998_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN1[20]),
    .B(_0085_),
    .X(_0491_)
);

sky130_fd_sc_hd__and2_4 _0999_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN7[20]),
    .B(_0197_),
    .X(_0492_)
);

sky130_fd_sc_hd__a21o_4 _1000_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN5[20]),
    .A2(_0241_),
    .B1(_0492_),
    .X(_0493_)
);

sky130_fd_sc_hd__and2_4 _1001_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN8[20]),
    .B(_0098_),
    .X(_0494_)
);

sky130_fd_sc_hd__a21o_4 _1002_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN2[20]),
    .A2(_0113_),
    .B1(_0494_),
    .X(_0495_)
);

sky130_fd_sc_hd__a21o_4 _1003_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN6[20]),
    .A2(_0090_),
    .B1(_0109_),
    .X(_0496_)
);

sky130_fd_sc_hd__and2_4 _1004_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(PAR_IN3[20]),
    .B(_0106_),
    .X(_0497_)
);

sky130_fd_sc_hd__a21o_4 _1005_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(PAR_IN4[20]),
    .A2(_0185_),
    .B1(_0497_),
    .X(_0498_)
);

sky130_fd_sc_hd__or4_4 _1006_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0493_),
    .B(_0495_),
    .C(_0496_),
    .D(_0498_),
    .X(_0499_)
);

sky130_fd_sc_hd__and3_4 _1007_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0122_),
    .B(_0491_),
    .C(_0499_),
    .X(_0500_)
);

sky130_fd_sc_hd__nor3_4 _1008_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0068_),
    .B(_0490_),
    .C(_0500_),
    .Y(_0501_)
);

sky130_fd_sc_hd__nor3_4 _1009_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0064_),
    .B(_0480_),
    .C(_0501_),
    .Y(_0502_)
);

sky130_fd_sc_hd__o21a_4 _1010_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0459_),
    .A2(_0502_),
    .B1(_0022_),
    .X(_0503_)
);

sky130_fd_sc_hd__nor3_4 _1011_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(COUNT[0]),
    .B(_0416_),
    .C(_0503_),
    .Y(_0504_)
);

sky130_fd_sc_hd__or4_4 _1012_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(SAMPLE_COUNT[3]),
    .B(COUNT[5]),
    .C(COMPLETE),
    .D(_0504_),
    .X(_0505_)
);

sky130_fd_sc_hd__nor2_4 _1013_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0328_),
    .B(_0505_),
    .Y(_0506_)
);

sky130_fd_sc_hd__a21o_4 _1014_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A1(_0040_),
    .A2(SERIAL_OUT),
    .B1(_0506_),
    .X(_0507_)
);

sky130_fd_sc_hd__and2_4 _1015_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(_0037_),
    .B(_0507_),
    .X(_0012_)
);

sky130_fd_sc_hd__dfrtp_4 _1016_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0012_),
    .Q(SERIAL_OUT),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1017_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0007_),
    .Q(INTERNAL_FINISH),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1018_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0000_),
    .Q(COMPLETE),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1019_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0001_),
    .Q(COUNT[0]),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1020_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0002_),
    .Q(COUNT[1]),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1021_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0003_),
    .Q(COUNT[2]),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1022_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0004_),
    .Q(COUNT[3]),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1023_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0005_),
    .Q(COUNT[4]),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1024_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0006_),
    .Q(COUNT[5]),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1025_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0008_),
    .Q(SAMPLE_COUNT[0]),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1026_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0009_),
    .Q(SAMPLE_COUNT[1]),
    .RESET_B(RESET),
    .CLK(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1027_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0010_),
    .Q(SAMPLE_COUNT[2]),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__dfrtp_4 _1028_ (
    .VGND(vgnd),
    .VPWR(vpwr),
    .D(_0011_),
    .Q(SAMPLE_COUNT[3]),
    .RESET_B(RESET),
    .CLK(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_96 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 PHY_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(CLK),
    .X(clknet_0_CLK)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_CLK),
    .X(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .A(clknet_0_CLK),
    .X(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_CLK_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1012__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COMPLETE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0562__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COMPLETE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0535__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COMPLETE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0528__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COMPLETE)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1011__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0835__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0560__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0558__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0516__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0923__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0833__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0560__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0517__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0921__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0832__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0740__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0515__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0570__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0513__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0889__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0868__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0855__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0628__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0509__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1012__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0580__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0557__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0521__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(COUNT[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0531__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(INTERNAL_FINISH)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0836__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0723__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0774__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0890__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0593__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0934__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0821__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0858__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0698__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0811__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0998__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0753__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0901__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0668__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0945__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0799__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0846__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0712__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0967__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0764__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0880__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0632__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0686__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0988__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0741__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0919__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0653__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0955__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0786__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN1[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0925__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0838__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0726__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0775__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0897__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0625__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0935__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0822__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0866__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0699__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0812__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0754__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0908__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0671__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0946__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0801__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0853__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0713__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0968__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0765__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0876__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0887__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0638__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0687__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0989__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0742__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0917__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0654__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0956__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0795__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN2[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0926__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0842__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0727__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0776__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0895__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0617__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0936__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0823__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0700__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0813__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1004__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0755__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0906__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0672__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0802__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0851__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0714__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0766__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0874__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0885__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0639__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0688__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0743__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0915__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0655__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0957__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0793__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN3[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0837__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0734__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0779__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0891__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0601__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0939__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0826__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0860__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0703__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0816__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1005__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0758__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0902__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0675__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0950__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0805__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0847__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0717__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0972__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0769__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0870__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0881__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0644__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0693__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0993__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0746__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0911__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0660__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0960__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0787__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN4[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0930__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0843__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0728__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0780__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0893__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0610__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0937__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0824__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0861__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0701__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0817__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1000__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0756__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0903__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0680__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0951__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0848__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0718__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0973__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0767__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0872__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0882__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0640__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0694__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0991__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0749__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0913__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0658__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0958__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN5[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0839__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0735__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0777__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0892__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0602__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0827__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0862__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0707__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0759__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0904__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0673__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0948__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0806__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0849__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0715__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0770__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0871__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0648__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0690__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0744__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0912__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0663__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0961__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0788__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN6[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0928__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0840__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0736__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0984__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0778__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0624__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0941__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0828__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0863__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0708__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0815__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0999__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0760__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0905__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0674__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0949__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0807__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0850__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0716__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0771__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0884__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0649__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0691__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0745__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0916__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0664__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN7[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0931__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0841__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[10])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0729__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[11])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0981__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[12])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0781__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[13])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0894__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[14])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0611__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[15])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[16])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0825__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[17])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[18])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0702__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[19])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0818__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1001__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[20])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0757__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[21])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[22])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0681__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[23])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[24])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0804__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[25])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0852__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[26])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0719__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[27])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0974__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[28])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0768__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[29])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0873__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0886__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[30])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0641__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[31])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0695__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0992__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[4])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0750__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[5])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0914__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[6])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0659__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[7])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0959__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[8])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0791__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(PAR_IN8[9])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0581__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(READY)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0532__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(READY)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1027__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1025__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1024__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1023__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1021__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1019__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1017__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__RESET_B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(RESET)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0598__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0537__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0508__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[0])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0544__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0542__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[1])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0603__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0594__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0585__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0551__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[2])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1012__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0587__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0541__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__0525__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SAMPLE_COUNT[3])
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(SERIAL_OUT)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0000_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1019__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0001_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0002_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1021__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0003_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0004_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1023__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0005_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1024__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0006_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1017__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0007_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1025__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0008_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0009_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1027__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0010_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0011_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0012_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0618__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0603__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0594__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0543__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0530__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0013_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0919__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0014_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0510__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0014_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0899__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0878__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0845__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0584__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0511__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0015_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0997__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0933__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0512__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0016_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0783__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0752__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0738__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0578__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0522__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0017_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0856__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0018_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0514__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0018_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0900__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0810__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0574__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0520__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0019_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0922__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0020_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0565__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0020_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0519__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0020_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0557__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0021_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0518__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0021_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0022_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0834__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0022_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0563__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0022_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0518__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0022_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0567__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0023_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0560__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0023_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0519__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0023_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0566__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0024_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0520__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0024_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0577__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0025_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0572__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0025_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0522__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0025_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0522__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0026_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0523__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0027_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0573__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0561__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0546__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0536__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0524__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0028_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0579__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0029_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0567__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0029_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0543__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0029_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0530__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0029_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0603__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0030_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0598__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0030_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0594__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0030_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0526__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0030_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0621__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0618__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0612__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0607__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0527__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0031_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0559__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0558__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0536__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0532__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0530__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0032_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0552__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0033_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0529__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0033_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0582__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0580__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0555__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0549__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0530__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0034_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0540__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0035_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0582__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0036_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0532__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0036_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0037_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0580__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0037_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0556__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0037_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0533__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0037_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0562__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0038_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0534__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0038_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0583__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0558__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0555__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0548__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0540__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0039_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0582__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0558__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0548__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0539__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0040_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0582__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0041_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0539__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0041_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0586__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0042_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0538__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0042_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0621__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0612__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0607__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0546__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0539__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0043_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0540__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0044_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0577__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0575__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0557__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0550__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0547__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0045_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0621__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0612__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0603__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0598__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0543__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0046_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0552__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0047_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0547__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0047_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0586__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0048_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0545__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0048_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0618__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0607__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0594__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0548__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0546__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0049_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0547__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0050_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0549__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0051_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0549__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0052_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0580__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0568__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0563__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0556__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0555__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0053_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0621__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0607__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0581__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0554__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0553__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0054_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0581__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0055_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0554__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0055_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0553__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0055_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0555__C1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0056_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0556__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0057_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0555__D1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0057_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0558__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0058_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0581__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0579__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0576__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0569__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0564__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0059_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0561__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0060_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0564__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0061_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0578__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0062_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0575__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0062_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0568__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0062_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0563__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0062_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0564__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0063_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0785__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0685__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0568__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0567__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0064_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0572__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0065_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0567__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0065_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0569__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0066_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0569__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0067_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0944__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0920__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0571__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0068_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0831__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0763__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0711__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0684__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0572__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0069_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0573__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0070_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0576__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0071_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0965__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0784__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0739__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0652__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0575__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0072_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0576__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0073_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0578__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0074_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0579__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0075_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0583__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0076_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0964__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0820__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0697__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0666__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0627__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0077_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0618__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0078_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0612__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0078_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0598__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0078_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0586__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0078_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0587__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0079_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0588__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0080_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0864__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0851__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0841__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0615__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0589__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0081_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0906__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0895__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0885__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0874__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0590__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0082_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0846__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0836__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0591__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0083_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0924__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0919__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0798__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0630__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0592__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0084_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0998__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0821__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0722__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0686__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0593__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0085_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0627__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0086_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0849__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0087_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0087_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0646__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0087_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0595__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0087_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0904__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0883__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0862__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0661__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0596__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0088_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0994__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0983__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0961__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0806__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0597__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0089_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0777__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0770__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0759__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0602__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0090_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0859__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0091_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0847__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0091_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0837__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0091_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0599__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0091_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0911__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0787__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0730__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0692__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0600__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0092_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0972__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0939__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0642__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0601__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0093_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0602__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0094_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0626__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0095_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0886__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0865__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0852__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0604__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0096_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0907__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0894__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0873__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0841__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0605__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0097_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0914__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0676__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0656__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0606__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0098_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0825__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0818__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0641__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0611__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0099_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0893__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0872__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0608__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0100_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0913__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0848__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0747__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0678__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0609__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0101_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0824__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0817__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0658__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0640__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0610__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0102_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0611__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0103_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0626__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0104_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0851__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0842__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0633__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0613__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0105_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1004__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0915__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0906__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0724__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0614__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0106_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0957__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0823__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0813__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0688__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0617__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0107_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0915__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0792__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0732__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0643__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0616__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0108_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1003__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0826__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0816__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0693__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0617__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0109_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0626__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0110_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0800__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0669__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0636__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0619__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0111_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0968__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0925__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0897__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0887__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0620__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0112_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0795__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0775__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0765__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0625__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0113_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0896__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0114_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0875__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0114_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0704__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0114_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0622__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0114_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0916__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0863__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0850__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0840__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0623__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0115_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0928__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0689__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0645__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0624__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0116_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0625__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0117_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0626__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0118_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0627__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0119_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0652__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0120_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0943__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0629__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0121_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0830__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0809__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0667__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0651__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0122_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0967__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0945__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0934__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0631__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0123_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0712__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0698__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0668__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0653__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0632__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0124_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0651__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0125_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0895__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0885__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0874__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0864__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0634__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0126_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0936__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0926__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0635__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0127_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0714__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0700__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0672__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0655__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0639__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0128_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0876__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0866__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0853__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0838__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0637__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0129_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0917__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0699__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0687__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0654__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0638__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0130_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0639__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0131_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0650__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0132_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0641__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0133_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0650__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0134_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0717__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0703__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0675__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0660__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0644__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0135_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0717__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0703__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0675__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0660__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0644__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0136_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0650__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0137_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0745__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0716__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0674__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0664__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0649__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0138_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0970__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0927__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0892__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0871__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0647__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0139_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0827__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0715__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0690__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0673__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0648__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0140_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0649__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0141_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0650__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0142_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0651__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0143_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0652__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0144_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0685__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0145_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0666__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0146_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0655__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0147_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0665__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0148_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0981__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0931__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0791__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0657__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0149_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0729__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0719__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0702__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0695__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0659__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0150_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0659__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0151_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0665__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0152_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0665__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0153_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0948__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0940__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0912__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0814__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0662__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0154_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0788__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0744__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0735__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0707__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0663__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0155_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0664__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0156_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0665__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0157_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0666__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0158_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0684__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0159_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0773__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0762__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0710__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0160_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0683__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0161_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0978__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0946__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0935__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0670__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0162_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0754__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0742__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0726__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0671__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0163_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0672__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0164_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0682__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0165_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0674__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0166_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0682__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0167_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0682__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0168_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0992__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0974__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0959__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0804__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0677__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0169_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0781__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0768__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0757__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0750__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0681__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0170_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0980__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0937__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0930__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0171_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0728__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0718__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0701__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0694__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0680__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0172_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0681__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0173_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0682__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0174_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0683__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0175_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0684__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0176_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0685__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0177_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0834__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0178_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0697__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0179_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0688__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0180_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0696__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0181_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0828__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0807__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0691__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0182_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0691__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0183_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0696__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0184_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1005__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0960__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0826__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0816__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0693__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0185_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0696__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0186_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0695__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0187_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0696__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0188_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0697__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0189_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0711__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0190_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0710__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0191_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0700__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0192_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0709__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0193_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0702__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0194_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0709__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0195_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0709__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0196_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0999__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0905__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0884__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0794__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0705__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0197_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0984__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0949__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0941__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0815__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0706__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0198_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0778__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0771__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0760__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0736__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0708__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0199_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0708__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0200_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0709__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0201_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0710__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0202_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0711__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0203_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0740__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0204_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0721__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0205_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0714__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0206_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0720__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0207_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0716__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0208_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0720__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0209_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0720__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0210_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0719__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0211_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0720__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0212_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0721__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0213_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0739__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0214_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0774__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0764__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0753__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0741__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0723__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0215_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0738__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0216_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0802__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0793__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0725__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0217_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0776__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0766__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0755__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0743__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0727__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0218_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0727__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0219_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0737__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0220_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0729__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0221_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0737__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0222_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0993__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0950__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0805__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0731__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0223_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0779__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0769__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0758__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0746__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0734__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0224_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0993__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0982__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0960__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0805__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0733__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0225_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0779__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0769__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0758__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0746__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0734__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0226_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0737__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0227_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0736__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0228_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0737__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0229_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0738__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0230_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0739__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0231_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0740__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0232_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0834__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0233_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0752__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0234_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0743__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0235_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0751__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0236_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0745__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0237_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0751__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0238_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0751__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0239_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0973__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0958__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0951__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0803__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0748__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0240_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1000__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0780__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0767__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0756__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0749__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0241_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0750__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0242_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0751__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0243_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0752__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0244_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0763__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0245_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0762__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0246_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0755__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0247_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0761__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0248_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0757__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0249_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0761__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0250_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0761__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0251_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0760__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0252_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0761__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0253_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0762__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0254_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0763__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0255_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0785__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0256_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0773__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0257_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0766__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0258_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0772__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0259_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0768__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0260_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0772__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0261_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0772__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0262_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0771__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0263_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0772__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0264_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0773__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0265_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0784__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0266_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0783__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0267_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0776__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0268_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0782__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0269_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0778__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0270_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0782__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0271_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0782__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0272_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0781__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0273_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0782__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0274_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0783__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0275_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0784__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0276_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0785__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0277_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0834__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0278_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0797__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0279_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0788__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0280_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0796__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0281_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0903__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0882__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0861__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0843__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0790__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0282_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0791__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0283_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0796__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0284_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0972__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0950__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0939__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0929__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0793__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0285_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0796__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0286_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0795__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0287_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0796__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0288_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0797__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0289_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0810__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0290_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0988__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0977__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0955__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0811__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0799__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0291_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0809__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0292_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0956__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0908__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0822__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0812__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0801__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0293_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0802__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0294_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0808__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0295_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0804__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0296_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0808__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0297_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0808__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0298_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0807__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0299_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0808__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0300_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0809__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0301_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0810__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0302_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0832__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0303_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0820__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0304_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0813__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0305_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0819__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0306_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0815__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0307_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0819__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0308_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0819__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0309_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0818__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0310_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0819__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0311_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0820__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0312_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0831__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0313_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0830__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0314_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0823__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0315_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0829__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0316_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0825__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0317_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0829__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0318_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0829__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0319_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0828__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0320_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0829__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0321_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0830__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0322_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0831__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0323_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0832__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0324_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0833__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0325_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0834__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0326_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0835__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0327_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0328_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0845__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0329_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0838__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0330_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0844__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0331_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0840__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0332_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0844__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0333_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0844__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0334_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0843__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0335_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0844__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0336_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0845__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0337_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0856__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0338_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0855__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0339_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0848__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0340_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0854__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0341_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0850__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0342_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0854__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0343_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0854__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0344_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0853__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0345_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0854__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0346_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0855__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0347_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0856__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0348_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0922__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0349_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0901__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0890__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0880__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0869__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0858__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0350_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0868__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0351_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0902__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0891__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0881__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0870__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0860__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0352_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0861__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0353_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0354_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0863__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0355_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0867__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0356_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0867__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0357_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0866__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0358_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0867__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0359_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0868__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0360_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0879__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0361_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0878__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0362_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0871__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0363_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0877__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0364_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0873__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0365_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0877__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0366_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0877__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0367_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0876__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0368_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0877__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0369_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0878__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0370_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0879__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0371_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0922__A3 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0372_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0889__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0373_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0882__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0374_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0888__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0375_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0884__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0376_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0888__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0377_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0888__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0378_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0887__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0379_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0888__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0380_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0889__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0381_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0900__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0382_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0899__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0383_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0892__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0384_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0898__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0385_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0894__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0386_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0898__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0387_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0898__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0388_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0897__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0389_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0898__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0390_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0899__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0391_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0900__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0392_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0922__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0393_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0910__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0394_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0903__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0395_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0909__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0396_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0905__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0397_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0909__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0398_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0909__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0399_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0908__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0400_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0909__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0401_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0910__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0402_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0921__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0403_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0912__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0404_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0918__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0405_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0914__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0406_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0918__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0407_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0918__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0408_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0917__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0409_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0918__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0410_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0920__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0411_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0920__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0412_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0921__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0413_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0922__B2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0414_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0923__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0415_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1011__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0416_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0933__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0417_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0926__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0418_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0419_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0928__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0420_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0421_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0422_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0931__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0423_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0932__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0424_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0933__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0425_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0944__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0426_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0943__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0427_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0936__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0428_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0942__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0429_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0938__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0430_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0942__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0431_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0942__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0432_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0941__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0433_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0942__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0434_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0943__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0435_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0944__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0436_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0437_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0438_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0947__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0439_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0440_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0949__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0441_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0442_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0443_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0952__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0444_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0953__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0445_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0954__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0446_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0965__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0447_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0964__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0448_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0957__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0449_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0450_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0959__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0451_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0452_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0453_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0962__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0454_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0963__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0455_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0964__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0456_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0965__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0457_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0966__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0458_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__A1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0459_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0976__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0460_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0969__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0461_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0462_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0971__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0463_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0464_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0465_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0974__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0466_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0975__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0467_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0976__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0468_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0987__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0469_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0470_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0979__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0471_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0472_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0981__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0473_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0474_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0985__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0475_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0984__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0476_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0985__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0477_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0986__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0478_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0987__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0479_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0480_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0997__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0481_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0990__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0482_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0483_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0992__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0484_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0485_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0486_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0995__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0487_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0996__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0488_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__0997__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0489_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0490_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0491_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1000__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0492_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0493_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1002__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0494_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0495_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0496_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1005__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0497_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1006__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0498_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1007__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0499_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1008__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0500_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1009__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0501_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1010__A2 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0502_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1011__C (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0503_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1012__D (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0504_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0505_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1014__B1 (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0506_)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1015__B (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(_0507_)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_CLK_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_CLK_A (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1017__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1018__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1020__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1023__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1024__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1027__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1028__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_0_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1016__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1019__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1021__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1022__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1025__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__diode_2 ANTENNA__1026__CLK (
    .VGND(vgnd),
    .VPWR(vpwr),
    .DIODE(clknet_1_1_0_CLK)
);

sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_0_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_0_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_0_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_0_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_0_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_0_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_1_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_1_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_1_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_1_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_1_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_1_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_1_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_2_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_2_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_2_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_2_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_2_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_2_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_2_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_2_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_3_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_3_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_3_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_3_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_3_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_3_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_3_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_3_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_3_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_4_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_4_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_4_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_4_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_4_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_4_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_4_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_5_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_5_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_5_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_5_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_5_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_5_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_5_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_5_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_6_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_6_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_6_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_6_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_6_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_6_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_6_315 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_7_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_7_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_7_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_7_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_7_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_8_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_8_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_8_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_8_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_8_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_8_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_8_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_8_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_9_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_9_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_9_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_9_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_9_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_9_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_9_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_10_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_10_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_10_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_10_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_10_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_10_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_10_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_11_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_11_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_11_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_11_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_11_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_11_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_11_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_11_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_11_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_12_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_12_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_12_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_12_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_12_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_12_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_12_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_13_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_13_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_13_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_13_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_13_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_13_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_14_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_14_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_14_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_14_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_14_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_14_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_14_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_15_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_15_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_15_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_15_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_15_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_15_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_15_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_15_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_16_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_16_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_16_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_16_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_265 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_16_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_16_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_16_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_17_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_17_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_17_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_17_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_17_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_17_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_17_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_18_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_18_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_18_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_18_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_18_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_18_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_18_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_18_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_19_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_19_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_19_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_19_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_19_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_19_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_19_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_19_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_19_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_19_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_10 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_20_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_20_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_255 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_20_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_20_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_20_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_20_309 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_20_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_21_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_96 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_21_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_21_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_21_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_21_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_21_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_22_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_22_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_22_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_22_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_22_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_22_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_22_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_22_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_23_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_23_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_23_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_23_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_23_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_23_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_23_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_23_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_124 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_139 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_143 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_24_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_24_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_24_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_24_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_24_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_24_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_24_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_25_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_25_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_25_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_25_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_25_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_25_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_25_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_25_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_25_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_25_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_26_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_26_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_26_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_26_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_26_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_26_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_26_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_27_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_27_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_27_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_27_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_27_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_27_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_27_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_27_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_28_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_28_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_28_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_28_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_28_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_28_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_28_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_29_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_29_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_29_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_29_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_29_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_29_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_29_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_30_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_30_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_30_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_30_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_30_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_30_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_30_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_214 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_31_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_31_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_31_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_31_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_31_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_32_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_189 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_209 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_32_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_269 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_32_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_284 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_32_298 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_32_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_32_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_32_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_33_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_33_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_216 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_33_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_33_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_33_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_33_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_33_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_33_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_126 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_34_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_34_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_251 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_34_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_34_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_34_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_34_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_34_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_50 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_171 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_35_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_35_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_253 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_35_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_35_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_35_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_35_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_35_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_35_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_36_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_45 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_36_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_191 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_36_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_36_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_36_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_36_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_36_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_36_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_36_312 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_36_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_33 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_37_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_89 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_130 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_134 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_37_148 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_37_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_37_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_37_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_37_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_37_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_37 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_65 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_38_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_183 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_38_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_38_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_38_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_38_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_38_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_38_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_38_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_38_305 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_38_317 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_25 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_121 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_39_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_157 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_39_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_39_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_39_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_39_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_39_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_39_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_39_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_39_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_12 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_40_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_40_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_88 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_144 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_40_185 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_40_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_223 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_40_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_246 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_40_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_40_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_40_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_40_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_41_79 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_41_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_140 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_41_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_41_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_41_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_286 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_41_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_41_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_41_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_41_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_14 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_18 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_42_36 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_83 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_90 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_42_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_42_146 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_152 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_42_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_42_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_226 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_42_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_42_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_42_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_42_299 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_42_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_8 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_24 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_54 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_43_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_111 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_115 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_43_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_175 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_43_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_43_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_43_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_262 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_277 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_289 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_43_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_43_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_43_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_43_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_47 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_44_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_129 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_141 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_44_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_44_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_252 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_44_272 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_44_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_44_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_44_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_45_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_13 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_26 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_48 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_60 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_45_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_98 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_45_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_45_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_153 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_161 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_170 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_174 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_190 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_194 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_201 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_239 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_243 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_45_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_278 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_282 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_288 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_301 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_45_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_45_314 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_45_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_41 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_46 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_58 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_73 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_77 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_46_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_103 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_107 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_119 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_46_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_46_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_179 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_46_197 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_229 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_234 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_46_248 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_260 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_264 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_46_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_46_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_46_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_46_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_46_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_17 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_29 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_34 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_51 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_55 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_59 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_67 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_71 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_85 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_91 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_95 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_99 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_109 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_47_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_163 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_167 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_193 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_205 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_220 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_238 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_47_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_281 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_47_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_47_300 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_47_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_47_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_22 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_30 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_38 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_42 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_82 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_86 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_128 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_136 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_166 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_178 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_200 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_204 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_48_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_213 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_225 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_228 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_232 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_235 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_48_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_257 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_48_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_287 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_48_291 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_48_296 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_48_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_48_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_7 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_21 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_31 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_66 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_70 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_74 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_78 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_49_92 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_104 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_108 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_112 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_116 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_138 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_142 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_150 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_155 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_159 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_49_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_182 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_188 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_192 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_196 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_199 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_203 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_217 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_221 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_233 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_237 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_250 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_49_266 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_275 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_279 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_283 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_49_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_303 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_49_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_49_310 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_49_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_50_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_19 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_52 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_69 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_81 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_97 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_101 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_105 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_113 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_117 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_122 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_133 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_160 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_164 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_176 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_208 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_212 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_219 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_231 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_244 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_247 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_50_256 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_50_268 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_50_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_50_293 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_50_297 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_50_308 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_50_316 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_9 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_23 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_51_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_35 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_39 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_53 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_62 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_76 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_100 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_114 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_123 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_127 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_131 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_145 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_151 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_165 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_169 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_173 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_177 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_181 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_184 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_202 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_222 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_227 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_51_240 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_259 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_263 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_267 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_271 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_285 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_51_290 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_51_294 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_51_302 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_51_306 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_51_318 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_11 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_20 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_28 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_40 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_52_43 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_49 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_57 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_61 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_64 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_68 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_72 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_80 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_84 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_93 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_102 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_110 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_120 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_132 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_135 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_52_147 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_154 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_158 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_162 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_172 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_186 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_206 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_210 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_215 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_224 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_3 FILLER_52_236 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_241 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_245 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_254 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_258 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_52_270 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_52_274 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_52_276 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_52_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_295 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_52_307 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_3 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_15 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_4 FILLER_53_27 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_32 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_44 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_56 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_63 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_75 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_87 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_94 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_106 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_118 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_125 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_137 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_149 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_156 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_168 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_180 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_53_187 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_1 FILLER_53_195 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_198 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__fill_2 FILLER_53_207 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_211 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_218 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_230 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_242 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_249 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_261 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_273 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_280 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_12 FILLER_53_292 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_6 FILLER_53_304 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

sky130_fd_sc_hd__decap_8 FILLER_53_311 (
    .VGND(vgnd),
    .VPWR(vpwr)
);

endmodule
