* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599603751605
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_599603751606
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599603751602
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_599603751609
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT Inverter2 GND VDD INP OUT
** N=32 EP=4 IP=31 FDC=28
M0 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2210 $Y=1130 $D=9
M1 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2640 $Y=1130 $D=9
M2 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3070 $Y=1130 $D=9
M3 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3500 $Y=1130 $D=9
M4 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3930 $Y=1130 $D=9
M5 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4360 $Y=1130 $D=9
M6 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4790 $Y=1130 $D=9
M7 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5220 $Y=1130 $D=9
M8 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5650 $Y=1130 $D=9
M9 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1985 $Y=7395 $D=79
M10 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2415 $Y=7395 $D=79
M11 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2845 $Y=7395 $D=79
M12 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3275 $Y=7395 $D=79
M13 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3705 $Y=7395 $D=79
M14 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4135 $Y=7395 $D=79
M15 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4565 $Y=7395 $D=79
M16 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4995 $Y=7395 $D=79
M17 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5425 $Y=7395 $D=79
M18 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5855 $Y=7395 $D=79
M19 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6285 $Y=7395 $D=79
M20 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6715 $Y=7395 $D=79
M21 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7145 $Y=7395 $D=79
M22 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7575 $Y=7395 $D=79
M23 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8005 $Y=7395 $D=79
M24 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8435 $Y=7395 $D=79
M25 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8865 $Y=7395 $D=79
M26 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=9295 $Y=7395 $D=79
X27 GND VDD Dpar a=48.4008 p=28.78 m=1 $[nwdiode] $X=860 $Y=7215 $D=191
.ENDS
***************************************
.SUBCKT Inv_Transmitter GND VDD VIN VOUT
** N=62 EP=4 IP=42 FDC=42
M0 4 VIN GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2860 $Y=1715 $D=9
M1 5 4 GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6295 $Y=1710 $D=9
M2 GND 4 5 GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6725 $Y=1710 $D=9
M3 5 4 GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7155 $Y=1710 $D=9
M4 4 VIN VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2635 $Y=7980 $D=79
M5 VDD VIN 4 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3065 $Y=7980 $D=79
M6 5 4 VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6070 $Y=7975 $D=79
M7 VDD 4 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6500 $Y=7975 $D=79
M8 5 4 VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6930 $Y=7975 $D=79
M9 VDD 4 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7360 $Y=7975 $D=79
M10 5 4 VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=7790 $Y=7975 $D=79
M11 VDD 4 5 VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=8220 $Y=7975 $D=79
X12 GND VDD Dpar a=11.524 p=15.02 m=1 $[nwdiode] $X=1510 $Y=7800 $D=191
X13 GND VDD Dpar a=20.7432 p=18.46 m=1 $[nwdiode] $X=4945 $Y=7795 $D=191
X30 GND VDD 5 VOUT Inverter2 $T=9575 575 0 0 $X=9830 $Y=925
.ENDS
***************************************
