VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

MACRO serializer_unit_cell_1
  CLASS BLOCK ;
  FOREIGN serializer_unit_cell_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 159.555 BY 170.275 ;
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END CLK
  PIN COMPLETE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END COMPLETE
  PIN COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END COUNT[0]
  PIN COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 155.555 160.520 159.555 161.120 ;
    END
  END COUNT[1]
  PIN COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 155.555 44.240 159.555 44.840 ;
    END
  END COUNT[2]
  PIN COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 166.275 73.050 170.275 ;
    END
  END COUNT[3]
  PIN COUNT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END COUNT[4]
  PIN COUNT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END COUNT[5]
  PIN INTERNAL_FINISH
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END INTERNAL_FINISH
  PIN PAR_IN1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 166.275 113.530 170.275 ;
    END
  END PAR_IN1[0]
  PIN PAR_IN1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 166.275 10.490 170.275 ;
    END
  END PAR_IN1[10]
  PIN PAR_IN1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 166.275 20.610 170.275 ;
    END
  END PAR_IN1[11]
  PIN PAR_IN1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END PAR_IN1[12]
  PIN PAR_IN1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END PAR_IN1[13]
  PIN PAR_IN1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END PAR_IN1[14]
  PIN PAR_IN1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 166.275 14.170 170.275 ;
    END
  END PAR_IN1[15]
  PIN PAR_IN1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 166.275 85.010 170.275 ;
    END
  END PAR_IN1[16]
  PIN PAR_IN1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END PAR_IN1[17]
  PIN PAR_IN1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END PAR_IN1[18]
  PIN PAR_IN1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END PAR_IN1[19]
  PIN PAR_IN1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END PAR_IN1[1]
  PIN PAR_IN1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END PAR_IN1[20]
  PIN PAR_IN1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END PAR_IN1[21]
  PIN PAR_IN1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.230 166.275 119.510 170.275 ;
    END
  END PAR_IN1[22]
  PIN PAR_IN1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 166.275 0.370 170.275 ;
    END
  END PAR_IN1[23]
  PIN PAR_IN1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END PAR_IN1[24]
  PIN PAR_IN1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.710 166.275 90.990 170.275 ;
    END
  END PAR_IN1[25]
  PIN PAR_IN1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END PAR_IN1[26]
  PIN PAR_IN1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 8.200 159.555 8.800 ;
    END
  END PAR_IN1[27]
  PIN PAR_IN1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 145.560 159.555 146.160 ;
    END
  END PAR_IN1[28]
  PIN PAR_IN1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END PAR_IN1[29]
  PIN PAR_IN1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END PAR_IN1[2]
  PIN PAR_IN1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END PAR_IN1[30]
  PIN PAR_IN1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END PAR_IN1[31]
  PIN PAR_IN1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END PAR_IN1[3]
  PIN PAR_IN1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 166.275 105.250 170.275 ;
    END
  END PAR_IN1[4]
  PIN PAR_IN1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 140.120 159.555 140.720 ;
    END
  END PAR_IN1[5]
  PIN PAR_IN1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END PAR_IN1[6]
  PIN PAR_IN1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END PAR_IN1[7]
  PIN PAR_IN1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END PAR_IN1[8]
  PIN PAR_IN1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END PAR_IN1[9]
  PIN PAR_IN2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 166.275 139.750 170.275 ;
    END
  END PAR_IN2[0]
  PIN PAR_IN2[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 112.920 159.555 113.520 ;
    END
  END PAR_IN2[10]
  PIN PAR_IN2[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END PAR_IN2[11]
  PIN PAR_IN2[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 166.275 54.650 170.275 ;
    END
  END PAR_IN2[12]
  PIN PAR_IN2[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END PAR_IN2[13]
  PIN PAR_IN2[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END PAR_IN2[14]
  PIN PAR_IN2[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 148.960 159.555 149.560 ;
    END
  END PAR_IN2[15]
  PIN PAR_IN2[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END PAR_IN2[16]
  PIN PAR_IN2[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END PAR_IN2[17]
  PIN PAR_IN2[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END PAR_IN2[18]
  PIN PAR_IN2[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 97.960 159.555 98.560 ;
    END
  END PAR_IN2[19]
  PIN PAR_IN2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END PAR_IN2[1]
  PIN PAR_IN2[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END PAR_IN2[20]
  PIN PAR_IN2[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END PAR_IN2[21]
  PIN PAR_IN2[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 163.920 159.555 164.520 ;
    END
  END PAR_IN2[22]
  PIN PAR_IN2[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 83.000 159.555 83.600 ;
    END
  END PAR_IN2[23]
  PIN PAR_IN2[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 166.275 50.510 170.275 ;
    END
  END PAR_IN2[24]
  PIN PAR_IN2[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END PAR_IN2[25]
  PIN PAR_IN2[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 166.275 109.390 170.275 ;
    END
  END PAR_IN2[26]
  PIN PAR_IN2[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 136.720 159.555 137.320 ;
    END
  END PAR_IN2[27]
  PIN PAR_IN2[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END PAR_IN2[28]
  PIN PAR_IN2[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 53.080 159.555 53.680 ;
    END
  END PAR_IN2[29]
  PIN PAR_IN2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 95.240 159.555 95.840 ;
    END
  END PAR_IN2[2]
  PIN PAR_IN2[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 166.275 8.190 170.275 ;
    END
  END PAR_IN2[30]
  PIN PAR_IN2[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END PAR_IN2[31]
  PIN PAR_IN2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 47.640 159.555 48.240 ;
    END
  END PAR_IN2[3]
  PIN PAR_IN2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END PAR_IN2[4]
  PIN PAR_IN2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END PAR_IN2[5]
  PIN PAR_IN2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 166.275 62.930 170.275 ;
    END
  END PAR_IN2[6]
  PIN PAR_IN2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END PAR_IN2[7]
  PIN PAR_IN2[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.910 166.275 123.190 170.275 ;
    END
  END PAR_IN2[8]
  PIN PAR_IN2[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END PAR_IN2[9]
  PIN PAR_IN3[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 17.720 159.555 18.320 ;
    END
  END PAR_IN3[0]
  PIN PAR_IN3[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END PAR_IN3[10]
  PIN PAR_IN3[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END PAR_IN3[11]
  PIN PAR_IN3[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END PAR_IN3[12]
  PIN PAR_IN3[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END PAR_IN3[13]
  PIN PAR_IN3[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END PAR_IN3[14]
  PIN PAR_IN3[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 134.000 159.555 134.600 ;
    END
  END PAR_IN3[15]
  PIN PAR_IN3[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 151.680 159.555 152.280 ;
    END
  END PAR_IN3[16]
  PIN PAR_IN3[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END PAR_IN3[17]
  PIN PAR_IN3[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 86.400 159.555 87.000 ;
    END
  END PAR_IN3[18]
  PIN PAR_IN3[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 166.275 77.190 170.275 ;
    END
  END PAR_IN3[19]
  PIN PAR_IN3[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END PAR_IN3[1]
  PIN PAR_IN3[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END PAR_IN3[20]
  PIN PAR_IN3[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 166.275 2.210 170.275 ;
    END
  END PAR_IN3[21]
  PIN PAR_IN3[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END PAR_IN3[22]
  PIN PAR_IN3[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 61.920 159.555 62.520 ;
    END
  END PAR_IN3[23]
  PIN PAR_IN3[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END PAR_IN3[24]
  PIN PAR_IN3[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END PAR_IN3[25]
  PIN PAR_IN3[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.310 166.275 141.590 170.275 ;
    END
  END PAR_IN3[26]
  PIN PAR_IN3[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END PAR_IN3[27]
  PIN PAR_IN3[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 155.080 159.555 155.680 ;
    END
  END PAR_IN3[28]
  PIN PAR_IN3[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END PAR_IN3[29]
  PIN PAR_IN3[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END PAR_IN3[2]
  PIN PAR_IN3[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END PAR_IN3[30]
  PIN PAR_IN3[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END PAR_IN3[31]
  PIN PAR_IN3[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 166.275 46.830 170.275 ;
    END
  END PAR_IN3[3]
  PIN PAR_IN3[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 166.275 44.530 170.275 ;
    END
  END PAR_IN3[4]
  PIN PAR_IN3[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 166.275 34.410 170.275 ;
    END
  END PAR_IN3[5]
  PIN PAR_IN3[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 2.760 159.555 3.360 ;
    END
  END PAR_IN3[6]
  PIN PAR_IN3[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END PAR_IN3[7]
  PIN PAR_IN3[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 166.275 12.330 170.275 ;
    END
  END PAR_IN3[8]
  PIN PAR_IN3[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 166.275 22.450 170.275 ;
    END
  END PAR_IN3[9]
  PIN PAR_IN4[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.150 166.275 143.430 170.275 ;
    END
  END PAR_IN4[0]
  PIN PAR_IN4[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 166.275 80.870 170.275 ;
    END
  END PAR_IN4[10]
  PIN PAR_IN4[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.030 166.275 133.310 170.275 ;
    END
  END PAR_IN4[11]
  PIN PAR_IN4[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END PAR_IN4[12]
  PIN PAR_IN4[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 89.120 159.555 89.720 ;
    END
  END PAR_IN4[13]
  PIN PAR_IN4[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 121.760 159.555 122.360 ;
    END
  END PAR_IN4[14]
  PIN PAR_IN4[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END PAR_IN4[15]
  PIN PAR_IN4[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 59.200 159.555 59.800 ;
    END
  END PAR_IN4[16]
  PIN PAR_IN4[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 50.360 159.555 50.960 ;
    END
  END PAR_IN4[17]
  PIN PAR_IN4[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 20.440 159.555 21.040 ;
    END
  END PAR_IN4[18]
  PIN PAR_IN4[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 166.275 40.850 170.275 ;
    END
  END PAR_IN4[19]
  PIN PAR_IN4[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 166.275 79.030 170.275 ;
    END
  END PAR_IN4[1]
  PIN PAR_IN4[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END PAR_IN4[20]
  PIN PAR_IN4[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END PAR_IN4[21]
  PIN PAR_IN4[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END PAR_IN4[22]
  PIN PAR_IN4[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.270 166.275 153.550 170.275 ;
    END
  END PAR_IN4[23]
  PIN PAR_IN4[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 166.275 93.290 170.275 ;
    END
  END PAR_IN4[24]
  PIN PAR_IN4[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 166.275 6.350 170.275 ;
    END
  END PAR_IN4[25]
  PIN PAR_IN4[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 166.275 52.810 170.275 ;
    END
  END PAR_IN4[26]
  PIN PAR_IN4[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END PAR_IN4[27]
  PIN PAR_IN4[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END PAR_IN4[28]
  PIN PAR_IN4[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END PAR_IN4[29]
  PIN PAR_IN4[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 74.160 159.555 74.760 ;
    END
  END PAR_IN4[2]
  PIN PAR_IN4[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 166.275 135.610 170.275 ;
    END
  END PAR_IN4[30]
  PIN PAR_IN4[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 166.275 115.370 170.275 ;
    END
  END PAR_IN4[31]
  PIN PAR_IN4[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 41.520 159.555 42.120 ;
    END
  END PAR_IN4[3]
  PIN PAR_IN4[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END PAR_IN4[4]
  PIN PAR_IN4[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END PAR_IN4[5]
  PIN PAR_IN4[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END PAR_IN4[6]
  PIN PAR_IN4[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 104.080 159.555 104.680 ;
    END
  END PAR_IN4[7]
  PIN PAR_IN4[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END PAR_IN4[8]
  PIN PAR_IN4[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.350 166.275 129.630 170.275 ;
    END
  END PAR_IN4[9]
  PIN PAR_IN5[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 166.275 64.770 170.275 ;
    END
  END PAR_IN5[0]
  PIN PAR_IN5[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END PAR_IN5[10]
  PIN PAR_IN5[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END PAR_IN5[11]
  PIN PAR_IN5[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END PAR_IN5[12]
  PIN PAR_IN5[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END PAR_IN5[13]
  PIN PAR_IN5[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 166.275 89.150 170.275 ;
    END
  END PAR_IN5[14]
  PIN PAR_IN5[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END PAR_IN5[15]
  PIN PAR_IN5[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END PAR_IN5[16]
  PIN PAR_IN5[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END PAR_IN5[17]
  PIN PAR_IN5[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END PAR_IN5[18]
  PIN PAR_IN5[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END PAR_IN5[19]
  PIN PAR_IN5[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END PAR_IN5[1]
  PIN PAR_IN5[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 166.275 58.790 170.275 ;
    END
  END PAR_IN5[20]
  PIN PAR_IN5[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END PAR_IN5[21]
  PIN PAR_IN5[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 166.275 60.630 170.275 ;
    END
  END PAR_IN5[22]
  PIN PAR_IN5[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 166.275 107.090 170.275 ;
    END
  END PAR_IN5[23]
  PIN PAR_IN5[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 166.275 159.530 170.275 ;
    END
  END PAR_IN5[24]
  PIN PAR_IN5[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 166.275 24.290 170.275 ;
    END
  END PAR_IN5[25]
  PIN PAR_IN5[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 110.200 159.555 110.800 ;
    END
  END PAR_IN5[26]
  PIN PAR_IN5[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END PAR_IN5[27]
  PIN PAR_IN5[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 76.880 159.555 77.480 ;
    END
  END PAR_IN5[28]
  PIN PAR_IN5[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END PAR_IN5[29]
  PIN PAR_IN5[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END PAR_IN5[2]
  PIN PAR_IN5[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 38.120 159.555 38.720 ;
    END
  END PAR_IN5[30]
  PIN PAR_IN5[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END PAR_IN5[31]
  PIN PAR_IN5[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 166.275 26.590 170.275 ;
    END
  END PAR_IN5[3]
  PIN PAR_IN5[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END PAR_IN5[4]
  PIN PAR_IN5[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 115.640 159.555 116.240 ;
    END
  END PAR_IN5[5]
  PIN PAR_IN5[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END PAR_IN5[6]
  PIN PAR_IN5[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 166.275 18.310 170.275 ;
    END
  END PAR_IN5[7]
  PIN PAR_IN5[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END PAR_IN5[8]
  PIN PAR_IN5[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END PAR_IN5[9]
  PIN PAR_IN6[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END PAR_IN6[0]
  PIN PAR_IN6[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END PAR_IN6[10]
  PIN PAR_IN6[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 65.320 159.555 65.920 ;
    END
  END PAR_IN6[11]
  PIN PAR_IN6[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 166.275 67.070 170.275 ;
    END
  END PAR_IN6[12]
  PIN PAR_IN6[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END PAR_IN6[13]
  PIN PAR_IN6[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END PAR_IN6[14]
  PIN PAR_IN6[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END PAR_IN6[15]
  PIN PAR_IN6[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END PAR_IN6[16]
  PIN PAR_IN6[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END PAR_IN6[17]
  PIN PAR_IN6[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.130 166.275 103.410 170.275 ;
    END
  END PAR_IN6[18]
  PIN PAR_IN6[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 166.275 48.670 170.275 ;
    END
  END PAR_IN6[19]
  PIN PAR_IN6[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 166.275 32.570 170.275 ;
    END
  END PAR_IN6[1]
  PIN PAR_IN6[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 130.600 159.555 131.200 ;
    END
  END PAR_IN6[20]
  PIN PAR_IN6[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 166.275 38.550 170.275 ;
    END
  END PAR_IN6[21]
  PIN PAR_IN6[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END PAR_IN6[22]
  PIN PAR_IN6[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.590 166.275 149.870 170.275 ;
    END
  END PAR_IN6[23]
  PIN PAR_IN6[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 56.480 159.555 57.080 ;
    END
  END PAR_IN6[24]
  PIN PAR_IN6[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END PAR_IN6[25]
  PIN PAR_IN6[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END PAR_IN6[26]
  PIN PAR_IN6[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END PAR_IN6[27]
  PIN PAR_IN6[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END PAR_IN6[28]
  PIN PAR_IN6[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END PAR_IN6[29]
  PIN PAR_IN6[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 91.840 159.555 92.440 ;
    END
  END PAR_IN6[2]
  PIN PAR_IN6[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 29.280 159.555 29.880 ;
    END
  END PAR_IN6[30]
  PIN PAR_IN6[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END PAR_IN6[31]
  PIN PAR_IN6[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END PAR_IN6[3]
  PIN PAR_IN6[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 166.275 127.330 170.275 ;
    END
  END PAR_IN6[4]
  PIN PAR_IN6[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 166.275 95.130 170.275 ;
    END
  END PAR_IN6[5]
  PIN PAR_IN6[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 142.840 159.555 143.440 ;
    END
  END PAR_IN6[6]
  PIN PAR_IN6[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 166.275 16.470 170.275 ;
    END
  END PAR_IN6[7]
  PIN PAR_IN6[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END PAR_IN6[8]
  PIN PAR_IN6[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.470 166.275 70.750 170.275 ;
    END
  END PAR_IN6[9]
  PIN PAR_IN7[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 157.800 159.555 158.400 ;
    END
  END PAR_IN7[0]
  PIN PAR_IN7[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.210 166.275 125.490 170.275 ;
    END
  END PAR_IN7[10]
  PIN PAR_IN7[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 166.275 157.690 170.275 ;
    END
  END PAR_IN7[11]
  PIN PAR_IN7[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 101.360 159.555 101.960 ;
    END
  END PAR_IN7[12]
  PIN PAR_IN7[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END PAR_IN7[13]
  PIN PAR_IN7[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END PAR_IN7[14]
  PIN PAR_IN7[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END PAR_IN7[15]
  PIN PAR_IN7[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END PAR_IN7[16]
  PIN PAR_IN7[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 5.480 159.555 6.080 ;
    END
  END PAR_IN7[17]
  PIN PAR_IN7[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 166.275 147.570 170.275 ;
    END
  END PAR_IN7[18]
  PIN PAR_IN7[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END PAR_IN7[19]
  PIN PAR_IN7[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END PAR_IN7[1]
  PIN PAR_IN7[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 11.600 159.555 12.200 ;
    END
  END PAR_IN7[20]
  PIN PAR_IN7[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END PAR_IN7[21]
  PIN PAR_IN7[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END PAR_IN7[22]
  PIN PAR_IN7[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 166.275 56.950 170.275 ;
    END
  END PAR_IN7[23]
  PIN PAR_IN7[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 166.275 131.470 170.275 ;
    END
  END PAR_IN7[24]
  PIN PAR_IN7[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 166.275 117.210 170.275 ;
    END
  END PAR_IN7[25]
  PIN PAR_IN7[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END PAR_IN7[26]
  PIN PAR_IN7[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 166.275 151.710 170.275 ;
    END
  END PAR_IN7[27]
  PIN PAR_IN7[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 166.275 86.850 170.275 ;
    END
  END PAR_IN7[28]
  PIN PAR_IN7[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END PAR_IN7[29]
  PIN PAR_IN7[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 166.640 159.555 167.240 ;
    END
  END PAR_IN7[2]
  PIN PAR_IN7[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END PAR_IN7[30]
  PIN PAR_IN7[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 68.040 159.555 68.640 ;
    END
  END PAR_IN7[31]
  PIN PAR_IN7[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 166.275 137.450 170.275 ;
    END
  END PAR_IN7[3]
  PIN PAR_IN7[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 166.275 42.690 170.275 ;
    END
  END PAR_IN7[4]
  PIN PAR_IN7[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 166.275 155.850 170.275 ;
    END
  END PAR_IN7[5]
  PIN PAR_IN7[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END PAR_IN7[6]
  PIN PAR_IN7[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 166.275 99.270 170.275 ;
    END
  END PAR_IN7[7]
  PIN PAR_IN7[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 166.275 36.710 170.275 ;
    END
  END PAR_IN7[8]
  PIN PAR_IN7[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.450 166.275 145.730 170.275 ;
    END
  END PAR_IN7[9]
  PIN PAR_IN8[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.070 166.275 121.350 170.275 ;
    END
  END PAR_IN8[0]
  PIN PAR_IN8[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END PAR_IN8[10]
  PIN PAR_IN8[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END PAR_IN8[11]
  PIN PAR_IN8[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END PAR_IN8[12]
  PIN PAR_IN8[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 166.275 28.430 170.275 ;
    END
  END PAR_IN8[13]
  PIN PAR_IN8[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END PAR_IN8[14]
  PIN PAR_IN8[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 127.880 159.555 128.480 ;
    END
  END PAR_IN8[15]
  PIN PAR_IN8[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END PAR_IN8[16]
  PIN PAR_IN8[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END PAR_IN8[17]
  PIN PAR_IN8[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 14.320 159.555 14.920 ;
    END
  END PAR_IN8[18]
  PIN PAR_IN8[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 166.275 111.230 170.275 ;
    END
  END PAR_IN8[19]
  PIN PAR_IN8[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 166.275 74.890 170.275 ;
    END
  END PAR_IN8[1]
  PIN PAR_IN8[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END PAR_IN8[20]
  PIN PAR_IN8[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END PAR_IN8[21]
  PIN PAR_IN8[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END PAR_IN8[22]
  PIN PAR_IN8[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END PAR_IN8[23]
  PIN PAR_IN8[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END PAR_IN8[24]
  PIN PAR_IN8[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 166.275 96.970 170.275 ;
    END
  END PAR_IN8[25]
  PIN PAR_IN8[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 119.040 159.555 119.640 ;
    END
  END PAR_IN8[26]
  PIN PAR_IN8[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 26.560 159.555 27.160 ;
    END
  END PAR_IN8[27]
  PIN PAR_IN8[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 71.440 159.555 72.040 ;
    END
  END PAR_IN8[28]
  PIN PAR_IN8[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 35.400 159.555 36.000 ;
    END
  END PAR_IN8[29]
  PIN PAR_IN8[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END PAR_IN8[2]
  PIN PAR_IN8[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 80.280 159.555 80.880 ;
    END
  END PAR_IN8[30]
  PIN PAR_IN8[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END PAR_IN8[31]
  PIN PAR_IN8[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 166.275 101.110 170.275 ;
    END
  END PAR_IN8[3]
  PIN PAR_IN8[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 32.680 159.555 33.280 ;
    END
  END PAR_IN8[4]
  PIN PAR_IN8[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 125.160 159.555 125.760 ;
    END
  END PAR_IN8[5]
  PIN PAR_IN8[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END PAR_IN8[6]
  PIN PAR_IN8[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END PAR_IN8[7]
  PIN PAR_IN8[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 166.275 83.170 170.275 ;
    END
  END PAR_IN8[8]
  PIN PAR_IN8[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 166.275 68.910 170.275 ;
    END
  END PAR_IN8[9]
  PIN READY
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END READY
  PIN RESET
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 155.555 106.800 159.555 107.400 ;
    END
  END RESET
  PIN SAMPLE_COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END SAMPLE_COUNT[0]
  PIN SAMPLE_COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END SAMPLE_COUNT[1]
  PIN SAMPLE_COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.770 166.275 4.050 170.275 ;
    END
  END SAMPLE_COUNT[2]
  PIN SAMPLE_COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 166.275 30.730 170.275 ;
    END
  END SAMPLE_COUNT[3]
  PIN SERIAL_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 155.555 23.160 159.555 23.760 ;
    END
  END SERIAL_OUT
  PIN VDD
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 153.640 28.090 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 153.640 104.680 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 0.145 0.085 153.640 166.855 ;
      LAYER met1 ;
        RECT 0.070 0.040 159.550 167.240 ;
      LAYER met2 ;
        RECT 0.650 165.995 1.650 167.270 ;
        RECT 2.490 165.995 3.490 167.270 ;
        RECT 4.330 165.995 5.790 167.270 ;
        RECT 6.630 165.995 7.630 167.270 ;
        RECT 8.470 165.995 9.930 167.270 ;
        RECT 10.770 165.995 11.770 167.270 ;
        RECT 12.610 165.995 13.610 167.270 ;
        RECT 14.450 165.995 15.910 167.270 ;
        RECT 16.750 165.995 17.750 167.270 ;
        RECT 18.590 165.995 20.050 167.270 ;
        RECT 20.890 165.995 21.890 167.270 ;
        RECT 22.730 165.995 23.730 167.270 ;
        RECT 24.570 165.995 26.030 167.270 ;
        RECT 26.870 165.995 27.870 167.270 ;
        RECT 28.710 165.995 30.170 167.270 ;
        RECT 31.010 165.995 32.010 167.270 ;
        RECT 32.850 165.995 33.850 167.270 ;
        RECT 34.690 165.995 36.150 167.270 ;
        RECT 36.990 165.995 37.990 167.270 ;
        RECT 38.830 165.995 40.290 167.270 ;
        RECT 41.130 165.995 42.130 167.270 ;
        RECT 42.970 165.995 43.970 167.270 ;
        RECT 44.810 165.995 46.270 167.270 ;
        RECT 47.110 165.995 48.110 167.270 ;
        RECT 48.950 165.995 49.950 167.270 ;
        RECT 50.790 165.995 52.250 167.270 ;
        RECT 53.090 165.995 54.090 167.270 ;
        RECT 54.930 165.995 56.390 167.270 ;
        RECT 57.230 165.995 58.230 167.270 ;
        RECT 59.070 165.995 60.070 167.270 ;
        RECT 60.910 165.995 62.370 167.270 ;
        RECT 63.210 165.995 64.210 167.270 ;
        RECT 65.050 165.995 66.510 167.270 ;
        RECT 67.350 165.995 68.350 167.270 ;
        RECT 69.190 165.995 70.190 167.270 ;
        RECT 71.030 165.995 72.490 167.270 ;
        RECT 73.330 165.995 74.330 167.270 ;
        RECT 75.170 165.995 76.630 167.270 ;
        RECT 77.470 165.995 78.470 167.270 ;
        RECT 79.310 165.995 80.310 167.270 ;
        RECT 81.150 165.995 82.610 167.270 ;
        RECT 83.450 165.995 84.450 167.270 ;
        RECT 85.290 165.995 86.290 167.270 ;
        RECT 87.130 165.995 88.590 167.270 ;
        RECT 89.430 165.995 90.430 167.270 ;
        RECT 91.270 165.995 92.730 167.270 ;
        RECT 93.570 165.995 94.570 167.270 ;
        RECT 95.410 165.995 96.410 167.270 ;
        RECT 97.250 165.995 98.710 167.270 ;
        RECT 99.550 165.995 100.550 167.270 ;
        RECT 101.390 165.995 102.850 167.270 ;
        RECT 103.690 165.995 104.690 167.270 ;
        RECT 105.530 165.995 106.530 167.270 ;
        RECT 107.370 165.995 108.830 167.270 ;
        RECT 109.670 165.995 110.670 167.270 ;
        RECT 111.510 165.995 112.970 167.270 ;
        RECT 113.810 165.995 114.810 167.270 ;
        RECT 115.650 165.995 116.650 167.270 ;
        RECT 117.490 165.995 118.950 167.270 ;
        RECT 119.790 165.995 120.790 167.270 ;
        RECT 121.630 165.995 122.630 167.270 ;
        RECT 123.470 165.995 124.930 167.270 ;
        RECT 125.770 165.995 126.770 167.270 ;
        RECT 127.610 165.995 129.070 167.270 ;
        RECT 129.910 165.995 130.910 167.270 ;
        RECT 131.750 165.995 132.750 167.270 ;
        RECT 133.590 165.995 135.050 167.270 ;
        RECT 135.890 165.995 136.890 167.270 ;
        RECT 137.730 165.995 139.190 167.270 ;
        RECT 140.030 165.995 141.030 167.270 ;
        RECT 141.870 165.995 142.870 167.270 ;
        RECT 143.710 165.995 145.170 167.270 ;
        RECT 146.010 165.995 147.010 167.270 ;
        RECT 147.850 165.995 149.310 167.270 ;
        RECT 150.150 165.995 151.150 167.270 ;
        RECT 151.990 165.995 152.990 167.270 ;
        RECT 153.830 165.995 155.290 167.270 ;
        RECT 156.130 165.995 157.130 167.270 ;
        RECT 157.970 165.995 158.970 167.270 ;
        RECT 0.090 4.280 159.250 165.995 ;
        RECT 0.650 0.010 1.650 4.280 ;
        RECT 2.490 0.010 3.490 4.280 ;
        RECT 4.330 0.010 5.790 4.280 ;
        RECT 6.630 0.010 7.630 4.280 ;
        RECT 8.470 0.010 9.470 4.280 ;
        RECT 10.310 0.010 11.770 4.280 ;
        RECT 12.610 0.010 13.610 4.280 ;
        RECT 14.450 0.010 15.910 4.280 ;
        RECT 16.750 0.010 17.750 4.280 ;
        RECT 18.590 0.010 19.590 4.280 ;
        RECT 20.430 0.010 21.890 4.280 ;
        RECT 22.730 0.010 23.730 4.280 ;
        RECT 24.570 0.010 26.030 4.280 ;
        RECT 26.870 0.010 27.870 4.280 ;
        RECT 28.710 0.010 29.710 4.280 ;
        RECT 30.550 0.010 32.010 4.280 ;
        RECT 32.850 0.010 33.850 4.280 ;
        RECT 34.690 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.990 4.280 ;
        RECT 38.830 0.010 39.830 4.280 ;
        RECT 40.670 0.010 42.130 4.280 ;
        RECT 42.970 0.010 43.970 4.280 ;
        RECT 44.810 0.010 45.810 4.280 ;
        RECT 46.650 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.950 4.280 ;
        RECT 50.790 0.010 52.250 4.280 ;
        RECT 53.090 0.010 54.090 4.280 ;
        RECT 54.930 0.010 55.930 4.280 ;
        RECT 56.770 0.010 58.230 4.280 ;
        RECT 59.070 0.010 60.070 4.280 ;
        RECT 60.910 0.010 62.370 4.280 ;
        RECT 63.210 0.010 64.210 4.280 ;
        RECT 65.050 0.010 66.050 4.280 ;
        RECT 66.890 0.010 68.350 4.280 ;
        RECT 69.190 0.010 70.190 4.280 ;
        RECT 71.030 0.010 72.490 4.280 ;
        RECT 73.330 0.010 74.330 4.280 ;
        RECT 75.170 0.010 76.170 4.280 ;
        RECT 77.010 0.010 78.470 4.280 ;
        RECT 79.310 0.010 80.310 4.280 ;
        RECT 81.150 0.010 82.150 4.280 ;
        RECT 82.990 0.010 84.450 4.280 ;
        RECT 85.290 0.010 86.290 4.280 ;
        RECT 87.130 0.010 88.590 4.280 ;
        RECT 89.430 0.010 90.430 4.280 ;
        RECT 91.270 0.010 92.270 4.280 ;
        RECT 93.110 0.010 94.570 4.280 ;
        RECT 95.410 0.010 96.410 4.280 ;
        RECT 97.250 0.010 98.710 4.280 ;
        RECT 99.550 0.010 100.550 4.280 ;
        RECT 101.390 0.010 102.390 4.280 ;
        RECT 103.230 0.010 104.690 4.280 ;
        RECT 105.530 0.010 106.530 4.280 ;
        RECT 107.370 0.010 108.830 4.280 ;
        RECT 109.670 0.010 110.670 4.280 ;
        RECT 111.510 0.010 112.510 4.280 ;
        RECT 113.350 0.010 114.810 4.280 ;
        RECT 115.650 0.010 116.650 4.280 ;
        RECT 117.490 0.010 118.490 4.280 ;
        RECT 119.330 0.010 120.790 4.280 ;
        RECT 121.630 0.010 122.630 4.280 ;
        RECT 123.470 0.010 124.930 4.280 ;
        RECT 125.770 0.010 126.770 4.280 ;
        RECT 127.610 0.010 128.610 4.280 ;
        RECT 129.450 0.010 130.910 4.280 ;
        RECT 131.750 0.010 132.750 4.280 ;
        RECT 133.590 0.010 135.050 4.280 ;
        RECT 135.890 0.010 136.890 4.280 ;
        RECT 137.730 0.010 138.730 4.280 ;
        RECT 139.570 0.010 141.030 4.280 ;
        RECT 141.870 0.010 142.870 4.280 ;
        RECT 143.710 0.010 145.170 4.280 ;
        RECT 146.010 0.010 147.010 4.280 ;
        RECT 147.850 0.010 148.850 4.280 ;
        RECT 149.690 0.010 151.150 4.280 ;
        RECT 151.990 0.010 152.990 4.280 ;
        RECT 153.830 0.010 155.290 4.280 ;
        RECT 156.130 0.010 157.130 4.280 ;
        RECT 157.970 0.010 158.970 4.280 ;
      LAYER met3 ;
        RECT 4.400 166.240 155.155 166.640 ;
        RECT 0.020 164.920 156.130 166.240 ;
        RECT 4.400 163.520 155.155 164.920 ;
        RECT 0.020 162.200 156.130 163.520 ;
        RECT 4.400 161.520 156.130 162.200 ;
        RECT 4.400 160.800 155.155 161.520 ;
        RECT 0.020 160.120 155.155 160.800 ;
        RECT 0.020 158.800 156.130 160.120 ;
        RECT 4.400 157.400 155.155 158.800 ;
        RECT 0.020 156.080 156.130 157.400 ;
        RECT 4.400 154.680 155.155 156.080 ;
        RECT 0.020 152.680 156.130 154.680 ;
        RECT 4.400 151.280 155.155 152.680 ;
        RECT 0.020 149.960 156.130 151.280 ;
        RECT 4.400 148.560 155.155 149.960 ;
        RECT 0.020 147.240 156.130 148.560 ;
        RECT 4.400 146.560 156.130 147.240 ;
        RECT 4.400 145.840 155.155 146.560 ;
        RECT 0.020 145.160 155.155 145.840 ;
        RECT 0.020 143.840 156.130 145.160 ;
        RECT 4.400 142.440 155.155 143.840 ;
        RECT 0.020 141.120 156.130 142.440 ;
        RECT 4.400 139.720 155.155 141.120 ;
        RECT 0.020 137.720 156.130 139.720 ;
        RECT 4.400 136.320 155.155 137.720 ;
        RECT 0.020 135.000 156.130 136.320 ;
        RECT 4.400 133.600 155.155 135.000 ;
        RECT 0.020 132.280 156.130 133.600 ;
        RECT 4.400 131.600 156.130 132.280 ;
        RECT 4.400 130.880 155.155 131.600 ;
        RECT 0.020 130.200 155.155 130.880 ;
        RECT 0.020 128.880 156.130 130.200 ;
        RECT 4.400 127.480 155.155 128.880 ;
        RECT 0.020 126.160 156.130 127.480 ;
        RECT 4.400 124.760 155.155 126.160 ;
        RECT 0.020 122.760 156.130 124.760 ;
        RECT 4.400 121.360 155.155 122.760 ;
        RECT 0.020 120.040 156.130 121.360 ;
        RECT 4.400 118.640 155.155 120.040 ;
        RECT 0.020 117.320 156.130 118.640 ;
        RECT 4.400 116.640 156.130 117.320 ;
        RECT 4.400 115.920 155.155 116.640 ;
        RECT 0.020 115.240 155.155 115.920 ;
        RECT 0.020 113.920 156.130 115.240 ;
        RECT 4.400 112.520 155.155 113.920 ;
        RECT 0.020 111.200 156.130 112.520 ;
        RECT 4.400 109.800 155.155 111.200 ;
        RECT 0.020 108.480 156.130 109.800 ;
        RECT 4.400 107.800 156.130 108.480 ;
        RECT 4.400 107.080 155.155 107.800 ;
        RECT 0.020 106.400 155.155 107.080 ;
        RECT 0.020 105.080 156.130 106.400 ;
        RECT 4.400 103.680 155.155 105.080 ;
        RECT 0.020 102.360 156.130 103.680 ;
        RECT 4.400 100.960 155.155 102.360 ;
        RECT 0.020 98.960 156.130 100.960 ;
        RECT 4.400 97.560 155.155 98.960 ;
        RECT 0.020 96.240 156.130 97.560 ;
        RECT 4.400 94.840 155.155 96.240 ;
        RECT 0.020 93.520 156.130 94.840 ;
        RECT 4.400 92.840 156.130 93.520 ;
        RECT 4.400 92.120 155.155 92.840 ;
        RECT 0.020 91.440 155.155 92.120 ;
        RECT 0.020 90.120 156.130 91.440 ;
        RECT 4.400 88.720 155.155 90.120 ;
        RECT 0.020 87.400 156.130 88.720 ;
        RECT 4.400 86.000 155.155 87.400 ;
        RECT 0.020 84.000 156.130 86.000 ;
        RECT 4.400 82.600 155.155 84.000 ;
        RECT 0.020 81.280 156.130 82.600 ;
        RECT 4.400 79.880 155.155 81.280 ;
        RECT 0.020 78.560 156.130 79.880 ;
        RECT 4.400 77.880 156.130 78.560 ;
        RECT 4.400 77.160 155.155 77.880 ;
        RECT 0.020 76.480 155.155 77.160 ;
        RECT 0.020 75.160 156.130 76.480 ;
        RECT 4.400 73.760 155.155 75.160 ;
        RECT 0.020 72.440 156.130 73.760 ;
        RECT 4.400 71.040 155.155 72.440 ;
        RECT 0.020 69.040 156.130 71.040 ;
        RECT 4.400 67.640 155.155 69.040 ;
        RECT 0.020 66.320 156.130 67.640 ;
        RECT 4.400 64.920 155.155 66.320 ;
        RECT 0.020 63.600 156.130 64.920 ;
        RECT 4.400 62.920 156.130 63.600 ;
        RECT 4.400 62.200 155.155 62.920 ;
        RECT 0.020 61.520 155.155 62.200 ;
        RECT 0.020 60.200 156.130 61.520 ;
        RECT 4.400 58.800 155.155 60.200 ;
        RECT 0.020 57.480 156.130 58.800 ;
        RECT 4.400 56.080 155.155 57.480 ;
        RECT 0.020 54.760 156.130 56.080 ;
        RECT 4.400 54.080 156.130 54.760 ;
        RECT 4.400 53.360 155.155 54.080 ;
        RECT 0.020 52.680 155.155 53.360 ;
        RECT 0.020 51.360 156.130 52.680 ;
        RECT 4.400 49.960 155.155 51.360 ;
        RECT 0.020 48.640 156.130 49.960 ;
        RECT 4.400 47.240 155.155 48.640 ;
        RECT 0.020 45.240 156.130 47.240 ;
        RECT 4.400 43.840 155.155 45.240 ;
        RECT 0.020 42.520 156.130 43.840 ;
        RECT 4.400 41.120 155.155 42.520 ;
        RECT 0.020 39.800 156.130 41.120 ;
        RECT 4.400 39.120 156.130 39.800 ;
        RECT 4.400 38.400 155.155 39.120 ;
        RECT 0.020 37.720 155.155 38.400 ;
        RECT 0.020 36.400 156.130 37.720 ;
        RECT 4.400 35.000 155.155 36.400 ;
        RECT 0.020 33.680 156.130 35.000 ;
        RECT 4.400 32.280 155.155 33.680 ;
        RECT 0.020 30.280 156.130 32.280 ;
        RECT 4.400 28.880 155.155 30.280 ;
        RECT 0.020 27.560 156.130 28.880 ;
        RECT 4.400 26.160 155.155 27.560 ;
        RECT 0.020 24.840 156.130 26.160 ;
        RECT 4.400 24.160 156.130 24.840 ;
        RECT 4.400 23.440 155.155 24.160 ;
        RECT 0.020 22.760 155.155 23.440 ;
        RECT 0.020 21.440 156.130 22.760 ;
        RECT 4.400 20.040 155.155 21.440 ;
        RECT 0.020 18.720 156.130 20.040 ;
        RECT 4.400 17.320 155.155 18.720 ;
        RECT 0.020 15.320 156.130 17.320 ;
        RECT 4.400 13.920 155.155 15.320 ;
        RECT 0.020 12.600 156.130 13.920 ;
        RECT 4.400 11.200 155.155 12.600 ;
        RECT 0.020 9.880 156.130 11.200 ;
        RECT 4.400 9.200 156.130 9.880 ;
        RECT 4.400 8.480 155.155 9.200 ;
        RECT 0.020 7.800 155.155 8.480 ;
        RECT 0.020 6.480 156.130 7.800 ;
        RECT 4.400 5.080 155.155 6.480 ;
        RECT 0.020 3.760 156.130 5.080 ;
        RECT 4.400 2.360 155.155 3.760 ;
        RECT 0.020 0.175 156.130 2.360 ;
      LAYER met4 ;
        RECT 0.295 1.535 156.105 158.265 ;
  END
END serializer_unit_cell_1
END LIBRARY

