* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_3 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=0.59 W=0.55 m=1 r=0.932203 a=0.3245 p=2.28 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=0.59 W=0.87 m=1 r=1.47458 a=0.5133 p=2.92 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 5440 1 0 $X=-190 $Y=2480
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=4 FDC=8
*.SEEDPROM
X0 1 2 ICV_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_1 $T=0 5440 0 0 $X=-190 $Y=5200
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=4 FDC=16
*.SEEDPROM
X0 1 2 ICV_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_2 $T=0 10880 0 0 $X=-190 $Y=10640
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.05 W=0.55 m=1 r=0.52381 a=0.5775 p=3.2 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.05 W=0.87 m=1 r=0.828571 a=0.9135 p=3.84 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_6 VNB VPB VGND VPWR
** N=14 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.97 W=0.55 m=1 r=0.279188 a=1.0835 p=5.04 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.97 W=0.87 m=1 r=0.441624 a=1.7139 p=5.68 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_8 VNB VPB VGND VPWR
** N=16 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=2.89 W=0.55 m=1 r=0.190311 a=1.5895 p=6.88 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=2.89 W=0.87 m=1 r=0.301038 a=2.5143 p=7.52 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_5 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 0 1 180 $X=3950 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_6 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=3680 0 0 0 $X=3490 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__diode_2 VNB DIODE
** N=9 EP=2 IP=0 FDC=1
*.SEEDPROM
D0 VNB DIODE ndiode AREA=0.4347 PJ=2.64 m=1 ahftempperim=2.64 $X=155 $Y=195 $D=167
.ENDS
***************************************
.SUBCKT ICV_7 1 3 4
** N=4 EP=3 IP=10 FDC=2
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 4 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_12 VNB VPB VGND VPWR
** N=18 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=4.73 W=0.55 m=1 r=0.116279 a=2.6015 p=10.56 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=4.73 W=0.87 m=1 r=0.183932 a=4.1151 p=11.2 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__buf_1 VNB VPB A VPWR X VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND A 7 VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 X 7 VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR A 7 VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 X 7 VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_10 1 3
** N=3 EP=2 IP=7 FDC=1
*.SEEDPROM
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3
** N=3 EP=3 IP=5 FDC=5
*.SEEDPROM
X0 1 2 ICV_5 $T=2300 0 0 0 $X=2110 $Y=-240
X1 1 3 ICV_10 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and2_4 VNB VPB A B VPWR X VGND
** N=38 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 9 A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=760 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1335 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1765 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2195 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2625 $Y=235 $D=9
M6 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M7 VPWR B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1335 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1765 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2195 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2625 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_12 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=3220 0 0 0 $X=3030 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21o_4 VNB VPB B1 A2 A1 VPWR X VGND
** N=55 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=850 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1280 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1710 $Y=235 $D=9
M4 9 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2675 $Y=235 $D=9
M5 VGND B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3095 $Y=235 $D=9
M6 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3555 $Y=235 $D=9
M7 9 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3935 $Y=235 $D=9
M8 12 A1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4355 $Y=235 $D=9
M9 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4775 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=850 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1280 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1710 $Y=1485 $D=89
M14 9 B1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2675 $Y=1485 $D=89
M15 10 B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3095 $Y=1485 $D=89
M16 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3515 $Y=1485 $D=89
M17 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3935 $Y=1485 $D=89
M18 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4355 $Y=1485 $D=89
M19 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4775 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_20 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4
** N=4 EP=4 IP=6 FDC=4
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_12 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=7
*.SEEDPROM
X0 1 2 3 2 4 1 sky130_fd_sc_hd__buf_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 ICV_16 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5 6 7
** N=7 EP=7 IP=13 FDC=21
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 6 7 2 4 1 sky130_fd_sc_hd__a21o_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=5
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 ICV_16 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=15
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 ICV_16 $T=4140 0 0 0 $X=3950 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_7 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=5
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 2 5 1 sky130_fd_sc_hd__buf_1 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=13
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__and2_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or4_4 VNB VPB D C B A VPWR X VGND
** N=46 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 10 D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND C 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=950 $Y=235 $D=9
M2 10 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1370 $Y=235 $D=9
M3 VGND A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1790 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2320 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2740 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3160 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M8 11 D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M9 12 C 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=950 $Y=1485 $D=88
M10 13 B 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1370 $Y=1485 $D=88
M11 VPWR A 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1790 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2320 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2740 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3160 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_7 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=23
*.SEEDPROM
X0 1 2 4 5 6 2 3 1 sky130_fd_sc_hd__a21o_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 7 ICV_31 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=23
*.SEEDPROM
X0 1 2 3 ICV_16 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 5 6 7 2 4 1 sky130_fd_sc_hd__a21o_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_35 1 3 4 5 6
** N=6 EP=5 IP=8 FDC=4
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 5 6 ICV_7 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_36 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_37 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_9 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_36 $T=5980 0 0 0 $X=5790 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_7 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=22
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 4 5 6 2 3 1 sky130_fd_sc_hd__a21o_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=22
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 2 5 1 sky130_fd_sc_hd__a21o_4 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_42 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_43 1 3 4
** N=4 EP=3 IP=6 FDC=2
*.SEEDPROM
X1 1 3 4 ICV_7 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_44 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X1 1 2 3 2 4 1 sky130_fd_sc_hd__buf_1 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=20
*.SEEDPROM
X1 1 2 4 5 6 2 3 1 sky130_fd_sc_hd__a21o_4 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_46 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_47 1 3
** N=3 EP=2 IP=7 FDC=1
*.SEEDPROM
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_48 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=11 FDC=23
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 5 6 7 8 9 ICV_23 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_50 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_51 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_4 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_52 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_53 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 ICV_18 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or2_4 VNB VPB B A VPWR X VGND
** N=37 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1740 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2580 $Y=235 $D=9
M6 9 B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=455 $Y=1485 $D=89
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2160 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_54 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and3_4 VNB VPB A B C VPWR X VGND
** N=43 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 10 A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=775 $Y=235 $D=9
M1 11 B 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=8
M2 VGND C 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1680 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2255 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2685 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3115 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3545 $Y=235 $D=9
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=775 $Y=1485 $D=89
M8 9 B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1750 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2255 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2685 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3115 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3545 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_55 1 2 3 4 5 6 7
** N=7 EP=7 IP=11 FDC=17
*.SEEDPROM
X0 1 2 3 ICV_16 $T=5060 0 0 0 $X=4870 $Y=-240
X1 1 2 4 5 6 2 7 1 sky130_fd_sc_hd__and3_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor3_4 VNB VPB A B C VPWR Y VGND
** N=63 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3775 $Y=235 $D=9
M9 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4195 $Y=235 $D=9
M10 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4615 $Y=235 $D=9
M11 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5035 $Y=235 $D=9
M12 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M13 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M14 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M15 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M16 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M17 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M18 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M19 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
M20 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3775 $Y=1485 $D=89
M21 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4195 $Y=1485 $D=89
M22 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4615 $Y=1485 $D=89
M23 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5035 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__inv_8 VNB VPB A VPWR Y VGND
** N=48 EP=6 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=560 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=980 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1400 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1820 $Y=235 $D=9
M4 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2240 $Y=235 $D=9
M5 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2660 $Y=235 $D=9
M6 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3080 $Y=235 $D=9
M7 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3500 $Y=235 $D=9
M8 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=560 $Y=1485 $D=89
M9 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=980 $Y=1485 $D=89
M10 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1400 $Y=1485 $D=89
M11 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1820 $Y=1485 $D=89
M12 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2240 $Y=1485 $D=89
M13 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2660 $Y=1485 $D=89
M14 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3080 $Y=1485 $D=89
M15 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3500 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o21a_4 VNB VPB B1 A1 A2 VPWR X VGND
** N=53 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 9 B1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2640 $Y=235 $D=9
M5 12 B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3070 $Y=235 $D=9
M6 VGND A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M7 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4090 $Y=235 $D=9
M8 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4520 $Y=235 $D=9
M9 12 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4950 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=720 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1150 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1580 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2010 $Y=1485 $D=89
M14 9 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2460 $Y=1485 $D=89
M15 VPWR B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2890 $Y=1485 $D=89
M16 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3660 $Y=1485 $D=89
M17 9 A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4090 $Y=1485 $D=89
M18 11 A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4520 $Y=1485 $D=89
M19 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4950 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or3_4 VNB VPB C B A VPWR X VGND
** N=49 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 VGND C 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 9 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2185 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2605 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3025 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3445 $Y=235 $D=9
M7 10 C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M8 11 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=88
M9 VPWR A 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2185 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2605 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3025 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3445 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4_4 VNB VPB A B C D VPWR X VGND
** N=44 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 11 A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 12 B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=790 $Y=235 $D=8
M2 13 C 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1275 $Y=235 $D=8
M3 VGND D 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1860 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2335 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2755 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3175 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3595 $Y=235 $D=9
M8 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M9 VPWR B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M10 10 C VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1275 $Y=1485 $D=89
M11 VPWR D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1855 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2335 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2755 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3175 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3595 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor2_4 VNB VPB A B VPWR Y VGND
** N=51 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M9 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M10 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M11 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M12 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M13 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M14 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M15 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dfrtp_4 VNB VPB CLK D RESET_B VPWR Q VGND
** N=88 EP=8 IP=0 FDC=34
*.SEEDPROM
M0 VGND CLK 9 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 10 9 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 15 D VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2090 $Y=235 $D=9
M3 12 9 15 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=2565 $Y=235 $D=9
M4 18 10 12 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=3045 $Y=235 $D=9
M5 19 11 18 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3875 $Y=235 $D=8
M6 VGND RESET_B 19 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4235 $Y=235 $D=9
M7 11 12 VGND VNB nshort L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=4895 $Y=235 $D=9
M8 14 10 11 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5390 $Y=235 $D=9
M9 20 9 14 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5935 $Y=235 $D=9
M10 VGND 13 20 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M11 21 RESET_B VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=235 $D=9
M12 13 14 21 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7615 $Y=235 $D=9
M13 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8555 $Y=235 $D=9
M14 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8975 $Y=235 $D=9
M15 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9395 $Y=235 $D=9
M16 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9815 $Y=235 $D=9
M17 VPWR CLK 9 VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M18 10 9 VPWR VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M19 15 D VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2150 $Y=2065 $D=89
M20 12 10 15 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2610 $Y=2065 $D=89
M21 16 9 12 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3105 $Y=2065 $D=89
M22 VPWR 11 16 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3805 $Y=2065 $D=89
M23 16 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4290 $Y=2065 $D=89
M24 11 12 VPWR VPB phighvt L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=5275 $Y=1645 $D=89
M25 14 9 11 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5770 $Y=2065 $D=89
M26 17 10 14 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6200 $Y=2065 $D=89
M27 VPWR 13 17 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6620 $Y=2065 $D=89
M28 13 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=2065 $D=89
M29 VPWR 14 13 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7580 $Y=2065 $D=89
M30 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8555 $Y=1485 $D=89
M31 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8975 $Y=1485 $D=89
M32 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9395 $Y=1485 $D=89
M33 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9815 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_1 VNB VPB A X VPWR VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND 7 X VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 7 A VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR 7 X VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 7 A VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21oi_4 VNB VPB B1 A2 A1 Y VPWR VGND
** N=57 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2590 $Y=235 $D=9
M6 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3020 $Y=235 $D=9
M7 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3450 $Y=235 $D=9
M8 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3880 $Y=235 $D=9
M9 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4310 $Y=235 $D=9
M10 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4740 $Y=235 $D=9
M11 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5170 $Y=235 $D=9
M12 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M13 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M14 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M15 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M16 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2150 $Y=1485 $D=89
M17 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2590 $Y=1485 $D=89
M18 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3020 $Y=1485 $D=89
M19 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3450 $Y=1485 $D=89
M20 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3880 $Y=1485 $D=89
M21 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4310 $Y=1485 $D=89
M22 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4740 $Y=1485 $D=89
M23 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nand2_4 VNB VPB B A VPWR Y VGND
** N=50 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND B 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 8 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 Y A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2915 $Y=235 $D=9
M7 8 A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3335 $Y=235 $D=9
M8 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M9 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M10 Y B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M11 VPWR B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M12 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M13 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M14 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2915 $Y=1485 $D=89
M15 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3335 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a2111oi_4 VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
** N=104 EP=10 IP=0 FDC=40
*.SEEDPROM
M0 Y D1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND D1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y D1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1265 $Y=235 $D=9
M3 VGND D1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1695 $Y=235 $D=9
M4 Y C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2205 $Y=235 $D=9
M5 VGND C1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2635 $Y=235 $D=9
M6 Y C1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3065 $Y=235 $D=9
M7 VGND C1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3495 $Y=235 $D=9
M8 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4035 $Y=235 $D=9
M9 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4465 $Y=235 $D=9
M10 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4895 $Y=235 $D=9
M11 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5325 $Y=235 $D=9
M12 Y A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6305 $Y=235 $D=9
M13 14 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6735 $Y=235 $D=9
M14 Y A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7165 $Y=235 $D=9
M15 14 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7595 $Y=235 $D=9
M16 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8120 $Y=235 $D=9
M17 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8550 $Y=235 $D=9
M18 VGND A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8980 $Y=235 $D=9
M19 14 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9410 $Y=235 $D=9
M20 Y D1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=405 $Y=1485 $D=89
M21 11 D1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M22 Y D1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1265 $Y=1485 $D=89
M23 11 D1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1695 $Y=1485 $D=89
M24 12 C1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2125 $Y=1485 $D=89
M25 11 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2555 $Y=1485 $D=89
M26 12 C1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2985 $Y=1485 $D=89
M27 11 C1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3415 $Y=1485 $D=89
M28 12 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4365 $Y=1485 $D=89
M29 13 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4795 $Y=1485 $D=89
M30 12 B1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5225 $Y=1485 $D=89
M31 13 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5655 $Y=1485 $D=89
M32 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6095 $Y=1485 $D=89
M33 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6525 $Y=1485 $D=89
M34 VPWR A1 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6955 $Y=1485 $D=89
M35 13 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7405 $Y=1485 $D=89
M36 VPWR A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7955 $Y=1485 $D=89
M37 13 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8385 $Y=1485 $D=89
M38 VPWR A2 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8905 $Y=1485 $D=89
M39 13 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9335 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_56 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT serializer_unit_cell_1 VSS VDD CLK PAR_IN7<29> PAR_IN1<23> SAMPLE_COUNT<2> PAR_IN7<13> PAR_IN6<13> PAR_IN4<12> RESET INTERNAL_FINISH PAR_IN6<29> PAR_IN2<1> PAR_IN5<12> PAR_IN4<25> READY PAR_IN3<1> PAR_IN4<4> PAR_IN8<12> PAR_IN2<25>
+ PAR_IN6<25> PAR_IN5<4> PAR_IN5<29> COMPLETE COUNT<4> PAR_IN5<15> PAR_IN6<8> PAR_IN8<7> PAR_IN5<7> PAR_IN3<12> COUNT<5> PAR_IN3<8> PAR_IN8<21> PAR_IN5<13> COUNT<1> PAR_IN1<24> COUNT<0> PAR_IN7<25> SAMPLE_COUNT<3> PAR_IN5<21>
+ PAR_IN7<8> PAR_IN3<25> PAR_IN4<8> PAR_IN5<8> PAR_IN8<13> PAR_IN1<12> PAR_IN5<25> PAR_IN1<26> SERIAL_OUT PAR_IN8<25> PAR_IN1<10> PAR_IN1<8> COUNT<3> PAR_IN8<8> PAR_IN4<20> PAR_IN3<20> PAR_IN3<4> PAR_IN7<4> COUNT<2> SAMPLE_COUNT<1>
+ SAMPLE_COUNT<0> PAR_IN6<26> PAR_IN8<4> PAR_IN2<12> PAR_IN6<21> PAR_IN6<4> PAR_IN2<5> PAR_IN2<4> PAR_IN3<9> PAR_IN7<26> PAR_IN3<5> PAR_IN3<13> PAR_IN1<9> PAR_IN2<24> PAR_IN2<31> PAR_IN2<7> PAR_IN1<18> PAR_IN4<5> PAR_IN3<31> PAR_IN1<2>
+ PAR_IN7<6> PAR_IN2<16> PAR_IN1<4> PAR_IN2<20> PAR_IN8<20> PAR_IN7<14> PAR_IN1<6> PAR_IN4<26> PAR_IN3<7> PAR_IN2<6> PAR_IN2<9> PAR_IN8<2> PAR_IN3<24> PAR_IN8<9> PAR_IN5<17> PAR_IN2<11> PAR_IN1<14> PAR_IN2<14> PAR_IN5<2> PAR_IN1<7>
+ PAR_IN8<10> PAR_IN3<11> PAR_IN5<20> PAR_IN1<13> PAR_IN3<29> PAR_IN1<31> PAR_IN6<9> PAR_IN6<0> PAR_IN3<21> PAR_IN1<20> PAR_IN8<29> PAR_IN8<6> PAR_IN2<21> PAR_IN8<14> PAR_IN1<25> PAR_IN4<29> PAR_IN8<17> PAR_IN1<16> PAR_IN8<22> PAR_IN1<15>
+ PAR_IN6<7> PAR_IN5<14> PAR_IN1<19> PAR_IN1<11> PAR_IN1<22> PAR_IN1<0> PAR_IN7<21> PAR_IN1<30> PAR_IN6<20> PAR_IN1<1> PAR_IN1<28> PAR_IN7<7> PAR_IN2<13> PAR_IN3<14> PAR_IN3<22> PAR_IN4<1> PAR_IN4<24> PAR_IN1<17> PAR_IN2<29> PAR_IN6<14>
+ PAR_IN6<15> PAR_IN1<27> PAR_IN3<6> PAR_IN2<22> PAR_IN7<15> PAR_IN5<3> PAR_IN4<13> PAR_IN4<15> PAR_IN8<1> PAR_IN2<15> PAR_IN6<5> PAR_IN4<21> PAR_IN3<17> PAR_IN8<15> PAR_IN8<3> PAR_IN1<29> PAR_IN1<3> PAR_IN7<5> PAR_IN1<5> PAR_IN3<15>
+ PAR_IN5<19> PAR_IN6<28> PAR_IN4<17> PAR_IN7<22> PAR_IN2<8> PAR_IN6<10> PAR_IN5<6> PAR_IN4<11> PAR_IN5<22> PAR_IN3<3> PAR_IN7<28> PAR_IN8<31> PAR_IN5<11> PAR_IN1<21> PAR_IN2<17> PAR_IN8<19> PAR_IN3<10> PAR_IN6<12> PAR_IN6<17> PAR_IN4<3>
+ PAR_IN4<10> PAR_IN8<24> PAR_IN6<22> PAR_IN5<0> PAR_IN5<23> PAR_IN6<3> PAR_IN8<11> PAR_IN5<10> PAR_IN7<10> PAR_IN5<27> PAR_IN5<26> PAR_IN6<1> PAR_IN5<31> PAR_IN5<1> PAR_IN7<3> PAR_IN4<19> PAR_IN2<26> PAR_IN7<17> PAR_IN3<30> PAR_IN5<9>
+ PAR_IN3<19> PAR_IN7<12> PAR_IN6<19> PAR_IN4<31> PAR_IN8<23> PAR_IN2<10> PAR_IN7<1> PAR_IN6<16> PAR_IN4<9> PAR_IN6<18> PAR_IN8<16> PAR_IN7<16> PAR_IN4<6> PAR_IN7<19> PAR_IN3<26> PAR_IN2<3> PAR_IN7<30> PAR_IN8<0> PAR_IN6<31> PAR_IN6<6>
+ PAR_IN3<2> PAR_IN2<30> PAR_IN8<27> PAR_IN7<24> PAR_IN7<31> PAR_IN2<19> PAR_IN6<30> PAR_IN7<18> PAR_IN5<16> PAR_IN7<23> PAR_IN3<18> PAR_IN5<18> PAR_IN7<11> PAR_IN4<28> PAR_IN6<27> PAR_IN8<18> PAR_IN7<0> PAR_IN3<27> PAR_IN2<18> PAR_IN3<16>
+ PAR_IN2<28> PAR_IN4<27> PAR_IN2<2> PAR_IN4<7> PAR_IN4<0> PAR_IN7<27> PAR_IN5<30> PAR_IN4<16> PAR_IN4<30> PAR_IN8<30> PAR_IN3<0> PAR_IN6<11> PAR_IN6<24> PAR_IN6<23> PAR_IN4<23> PAR_IN7<9> PAR_IN4<14> PAR_IN5<5> PAR_IN2<0> PAR_IN6<2>
+ PAR_IN8<5> PAR_IN3<28> PAR_IN7<20> PAR_IN3<23> PAR_IN8<28> PAR_IN7<2> PAR_IN8<26> PAR_IN4<22> PAR_IN2<27> PAR_IN4<18> PAR_IN4<2> PAR_IN5<28> PAR_IN5<24> PAR_IN2<23>
** N=1125 EP=274 IP=7642 FDC=11404
M0 26 3 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=17040 $Y=51915 $D=9
M1 VSS 3 26 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=17460 $Y=51915 $D=9
M2 26 3 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=17880 $Y=51915 $D=9
M3 VSS 3 26 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=18300 $Y=51915 $D=9
M4 3 4 40 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=19240 $Y=51915 $D=9
M5 40 5 3 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=19660 $Y=51915 $D=9
M6 3 5 40 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=20080 $Y=51915 $D=9
M7 40 4 3 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=20500 $Y=51915 $D=9
M8 VSS 6 40 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=21000 $Y=51915 $D=9
M9 40 7 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=21420 $Y=51915 $D=9
M10 9 CLK VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=21560 $Y=67345 $D=9
M11 VSS 7 40 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=21840 $Y=51915 $D=9
M12 VSS CLK 9 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=21990 $Y=67345 $D=9
M13 40 6 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=22260 $Y=51915 $D=9
M14 9 CLK VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=22420 $Y=67345 $D=9
M15 VSS CLK 9 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=22850 $Y=67345 $D=9
M16 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=23280 $Y=67345 $D=9
M17 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=23710 $Y=67345 $D=9
M18 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=24140 $Y=67345 $D=9
M19 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=24570 $Y=67345 $D=9
M20 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=25000 $Y=67345 $D=9
M21 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=25430 $Y=67345 $D=9
M22 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=25860 $Y=67345 $D=9
M23 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=26290 $Y=67345 $D=9
M24 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=26715 $Y=67345 $D=9
M25 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=27145 $Y=67345 $D=9
M26 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=27575 $Y=67345 $D=9
M27 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=28005 $Y=67345 $D=9
M28 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=28435 $Y=67345 $D=9
M29 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=28865 $Y=67345 $D=9
M30 29 9 VSS VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=29295 $Y=67345 $D=9
M31 VSS 9 29 VSS nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=29725 $Y=67345 $D=9
M32 30 10 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=35750 $Y=89995 $D=9
M33 VSS 10 30 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=36180 $Y=89995 $D=9
M34 30 10 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=36610 $Y=89995 $D=9
M35 VSS 10 30 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=37055 $Y=89995 $D=9
M36 10 11 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=37490 $Y=89995 $D=9
M37 VSS 12 10 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=37960 $Y=89995 $D=9
M38 10 12 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=38445 $Y=89995 $D=9
M39 VSS 11 10 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=38985 $Y=89995 $D=9
M40 41 13 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=39565 $Y=89995 $D=9
M41 10 14 41 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=39995 $Y=89995 $D=9
M42 42 14 10 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=40425 $Y=89995 $D=9
M43 VSS 13 42 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=40855 $Y=89995 $D=9
M44 34 15 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=56055 $Y=94315 $D=9
M45 VSS 15 34 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=56475 $Y=94315 $D=9
M46 34 15 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=56895 $Y=94315 $D=9
M47 VSS 15 34 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=57315 $Y=94315 $D=9
M48 43 16 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=57735 $Y=94315 $D=9
M49 VSS 16 43 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=58155 $Y=94315 $D=9
M50 43 17 44 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=59095 $Y=94315 $D=9
M51 44 17 43 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=59515 $Y=94315 $D=9
M52 15 18 44 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=59935 $Y=94315 $D=9
M53 44 18 15 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=60355 $Y=94315 $D=9
M54 15 19 45 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=61630 $Y=94315 $D=9
M55 45 19 15 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=62050 $Y=94315 $D=9
M56 VSS 20 45 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=62515 $Y=94315 $D=9
M57 45 20 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=62935 $Y=94315 $D=9
M58 37 21 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=68935 $Y=79115 $D=9
M59 46 21 37 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=69355 $Y=79115 $D=9
M60 37 21 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=69775 $Y=79115 $D=9
M61 46 21 37 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=70195 $Y=79115 $D=9
M62 37 22 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=70630 $Y=79115 $D=9
M63 46 22 37 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=71050 $Y=79115 $D=9
M64 37 22 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=71470 $Y=79115 $D=9
M65 46 22 37 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=71890 $Y=79115 $D=9
M66 VSS 23 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=72310 $Y=79115 $D=9
M67 46 23 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=72730 $Y=79115 $D=9
M68 VSS 23 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=73150 $Y=79115 $D=9
M69 46 23 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=73730 $Y=79115 $D=9
M70 VSS 24 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=74510 $Y=79115 $D=9
M71 46 24 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=74930 $Y=79115 $D=9
M72 VSS 24 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=75350 $Y=79115 $D=9
M73 46 24 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=75770 $Y=79115 $D=9
M74 VSS 25 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=76710 $Y=79115 $D=9
M75 46 25 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=77130 $Y=79115 $D=9
M76 VSS 25 46 VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=77550 $Y=79115 $D=9
M77 46 25 VSS VSS nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=78065 $Y=79115 $D=9
M78 26 3 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=17040 $Y=53165 $D=89
M79 VDD 3 26 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=17460 $Y=53165 $D=89
M80 26 3 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=17880 $Y=53165 $D=89
M81 VDD 3 26 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=18300 $Y=53165 $D=89
M82 27 4 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=19240 $Y=53165 $D=89
M83 3 5 27 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=19660 $Y=53165 $D=89
M84 27 5 3 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=20080 $Y=53165 $D=89
M85 VDD 4 27 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=20500 $Y=53165 $D=89
M86 28 6 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=21000 $Y=53165 $D=89
M87 3 7 28 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=21420 $Y=53165 $D=89
M88 9 CLK VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=21560 $Y=65515 $D=89
M89 28 7 3 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=21840 $Y=53165 $D=89
M90 VDD CLK 9 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=21990 $Y=65515 $D=89
M91 VDD 6 28 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=22260 $Y=53165 $D=89
M92 9 CLK VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=22420 $Y=65515 $D=89
M93 VDD CLK 9 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=22850 $Y=65515 $D=89
M94 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=23280 $Y=65515 $D=89
M95 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=23710 $Y=65515 $D=89
M96 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=24140 $Y=65515 $D=89
M97 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=24570 $Y=65515 $D=89
M98 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=25000 $Y=65515 $D=89
M99 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=25430 $Y=65515 $D=89
M100 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=25860 $Y=65515 $D=89
M101 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=26290 $Y=65515 $D=89
M102 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=26715 $Y=65515 $D=89
M103 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=27145 $Y=65515 $D=89
M104 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=27575 $Y=65515 $D=89
M105 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=28005 $Y=65515 $D=89
M106 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=28435 $Y=65515 $D=89
M107 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=28865 $Y=65515 $D=89
M108 29 9 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=29295 $Y=65515 $D=89
M109 VDD 9 29 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=29725 $Y=65515 $D=89
M110 30 10 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=35355 $Y=91245 $D=89
M111 VDD 10 30 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=35785 $Y=91245 $D=89
M112 30 10 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=36215 $Y=91245 $D=89
M113 VDD 10 30 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=36645 $Y=91245 $D=89
M114 32 11 31 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=37585 $Y=91245 $D=89
M115 10 12 32 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=38015 $Y=91245 $D=89
M116 33 12 10 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=38445 $Y=91245 $D=89
M117 31 11 33 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=38915 $Y=91245 $D=89
M118 VDD 13 31 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=39455 $Y=91245 $D=89
M119 31 14 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=39995 $Y=91245 $D=89
M120 VDD 14 31 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=40425 $Y=91245 $D=89
M121 31 13 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=40855 $Y=91245 $D=89
M122 34 15 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=56055 $Y=92715 $D=89
M123 VDD 15 34 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=56475 $Y=92715 $D=89
M124 34 15 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=56895 $Y=92715 $D=89
M125 VDD 15 34 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=57315 $Y=92715 $D=89
M126 35 16 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=57735 $Y=92715 $D=89
M127 VDD 16 35 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=58155 $Y=92715 $D=89
M128 VDD 17 35 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=59095 $Y=92715 $D=89
M129 35 17 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=59515 $Y=92715 $D=89
M130 VDD 18 35 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=59935 $Y=92715 $D=89
M131 35 18 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=60355 $Y=92715 $D=89
M132 15 19 35 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=61675 $Y=92715 $D=89
M133 35 19 15 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=62095 $Y=92715 $D=89
M134 15 20 35 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=62515 $Y=92715 $D=89
M135 35 20 15 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=62935 $Y=92715 $D=89
M136 37 21 36 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=68935 $Y=80365 $D=89
M137 36 21 37 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=69355 $Y=80365 $D=89
M138 37 21 36 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=69775 $Y=80365 $D=89
M139 36 21 37 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=70195 $Y=80365 $D=89
M140 VDD 22 36 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=70630 $Y=80365 $D=89
M141 36 22 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=71050 $Y=80365 $D=89
M142 VDD 22 36 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=71470 $Y=80365 $D=89
M143 36 22 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=71890 $Y=80365 $D=89
M144 37 23 38 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=72830 $Y=80365 $D=89
M145 38 23 37 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=73250 $Y=80365 $D=89
M146 37 23 38 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=73670 $Y=80365 $D=89
M147 38 23 37 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=74090 $Y=80365 $D=89
M148 39 24 38 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=74510 $Y=80365 $D=89
M149 38 24 39 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=74930 $Y=80365 $D=89
M150 39 24 38 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=75350 $Y=80365 $D=89
M151 38 24 39 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=75770 $Y=80365 $D=89
M152 39 25 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=76710 $Y=80365 $D=89
M153 VDD 25 39 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=77130 $Y=80365 $D=89
M154 39 25 VDD VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=77550 $Y=80365 $D=89
M155 VDD 25 39 VDD phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=78065 $Y=80365 $D=89
X156 VSS VDD Dpar a=238.342 p=300.21 m=1 $[nwdiode] $X=5330 $Y=10690 $D=191
X157 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=14905 $D=191
X158 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=20345 $D=191
X159 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=25785 $D=191
X160 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=31225 $D=191
X161 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=36665 $D=191
X162 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=42105 $D=191
X163 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=47545 $D=191
X164 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=52985 $D=191
X165 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=58425 $D=191
X166 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=63865 $D=191
X167 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=69305 $D=191
X168 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=74745 $D=191
X169 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=80185 $D=191
X170 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=85625 $D=191
X171 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=91065 $D=191
X172 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=96505 $D=191
X173 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=101945 $D=191
X174 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=107385 $D=191
X175 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=112825 $D=191
X176 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=118265 $D=191
X177 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=123705 $D=191
X178 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=129145 $D=191
X179 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=134585 $D=191
X180 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=140025 $D=191
X181 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=145465 $D=191
X182 VSS VDD Dpar a=420.255 p=302.66 m=1 $[nwdiode] $X=5330 $Y=150905 $D=191
X183 VSS VDD Dpar a=238.342 p=300.21 m=1 $[nwdiode] $X=5330 $Y=156345 $D=191
X184 806 VDD Probe probetype=1 $[VDD] $X=79578 $Y=27288 $D=314
X185 807 VSS Probe probetype=1 $[VSS] $X=79578 $Y=103878 $D=314
X186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 13600 1 0 $X=5330 $Y=10640
X187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 57120 1 0 $X=5330 $Y=54160
X188 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 116960 0 0 $X=5330 $Y=116720
X189 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=5520 155040 0 0 $X=5330 $Y=154800
X190 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=26680 138720 1 0 $X=26490 $Y=135760
X191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=32200 35360 0 0 $X=32010 $Y=35120
X192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=32660 13600 1 0 $X=32470 $Y=10640
X193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=48300 73440 1 0 $X=48110 $Y=70480
X194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=48300 78880 1 0 $X=48110 $Y=75920
X195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=55660 19040 1 0 $X=55470 $Y=16080
X196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=55660 106080 0 0 $X=55470 $Y=105840
X197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=59800 68000 1 0 $X=59610 $Y=65040
X198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=60260 95200 0 0 $X=60070 $Y=94960
X199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=62560 29920 1 0 $X=62370 $Y=26960
X200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=67160 51680 0 0 $X=66970 $Y=51440
X201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=76360 144160 1 0 $X=76170 $Y=141200
X202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=76360 149600 1 0 $X=76170 $Y=146640
X203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=80040 89760 1 0 $X=79850 $Y=86800
X204 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=80040 155040 1 0 $X=79850 $Y=152080
X205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=82340 122400 1 0 $X=82150 $Y=119440
X206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=94300 40800 1 0 $X=94110 $Y=37840
X207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=103500 19040 0 0 $X=103310 $Y=18800
X208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=115460 78880 1 0 $X=115270 $Y=75920
X209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=116380 84320 1 0 $X=116190 $Y=81360
X210 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=122360 13600 0 0 $X=122170 $Y=13360
X211 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=137540 89760 0 0 $X=137350 $Y=89520
X212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=142140 19040 1 0 $X=141950 $Y=16080
X213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=144440 84320 0 0 $X=144250 $Y=84080
X214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=150880 57120 1 0 $X=150690 $Y=54160
X215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 13600 0 180 $X=152070 $Y=10640
X216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 19040 0 180 $X=152070 $Y=16080
X217 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 24480 0 180 $X=152070 $Y=21520
X218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 35360 0 180 $X=152070 $Y=32400
X219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 51680 0 180 $X=152070 $Y=48720
X220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 57120 0 180 $X=152070 $Y=54160
X221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 62560 0 180 $X=152070 $Y=59600
X222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 73440 1 180 $X=152070 $Y=73200
X223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 89760 0 180 $X=152070 $Y=86800
X224 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 149600 0 180 $X=152070 $Y=146640
X225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3 $T=153640 155040 1 180 $X=152070 $Y=154800
X226 VSS VDD ICV_1 $T=5520 46240 0 0 $X=5330 $Y=46000
X227 VSS VDD ICV_1 $T=5520 100640 0 0 $X=5330 $Y=100400
X228 VSS VDD ICV_1 $T=5520 111520 0 0 $X=5330 $Y=111280
X229 VSS VDD ICV_1 $T=104420 24480 0 0 $X=104230 $Y=24240
X230 VSS VDD ICV_1 $T=153640 24480 1 180 $X=152070 $Y=24240
X231 VSS VDD ICV_1 $T=153640 78880 1 180 $X=152070 $Y=78640
X232 VSS VDD ICV_1 $T=153640 149600 1 180 $X=152070 $Y=149360
X233 VSS VDD ICV_2 $T=5520 35360 0 0 $X=5330 $Y=35120
X234 VSS VDD ICV_2 $T=153640 35360 1 180 $X=152070 $Y=35120
X235 VSS VDD ICV_2 $T=153640 62560 1 180 $X=152070 $Y=62320
X236 VSS VDD ICV_2 $T=153640 133280 1 180 $X=152070 $Y=133040
X237 VSS VDD ICV_3 $T=5520 13600 0 0 $X=5330 $Y=13360
X238 VSS VDD ICV_3 $T=5520 57120 0 0 $X=5330 $Y=56880
X239 VSS VDD ICV_3 $T=5520 78880 0 0 $X=5330 $Y=78640
X240 VSS VDD ICV_3 $T=5520 133280 0 0 $X=5330 $Y=133040
X241 VSS VDD ICV_3 $T=153640 89760 1 180 $X=152070 $Y=89520
X242 VSS VDD ICV_3 $T=153640 111520 1 180 $X=152070 $Y=111280
X243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=6900 40800 0 0 $X=6710 $Y=40560
X244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=12420 62560 0 0 $X=12230 $Y=62320
X245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=14260 51680 1 0 $X=14070 $Y=48720
X246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=16560 127840 0 0 $X=16370 $Y=127600
X247 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=18860 40800 0 0 $X=18670 $Y=40560
X248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=20240 40800 1 0 $X=20050 $Y=37840
X249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=23920 35360 0 0 $X=23730 $Y=35120
X250 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=28060 78880 0 0 $X=27870 $Y=78640
X251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=33580 116960 1 0 $X=33390 $Y=114000
X252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=40480 144160 1 0 $X=40290 $Y=141200
X253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=44620 138720 0 0 $X=44430 $Y=138480
X254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=53820 133280 1 0 $X=53630 $Y=130320
X255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=62100 127840 0 0 $X=61910 $Y=127600
X256 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=90160 95200 0 0 $X=89970 $Y=94960
X257 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=104420 35360 1 0 $X=104230 $Y=32400
X258 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=107180 144160 1 0 $X=106990 $Y=141200
X259 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=107640 111520 1 0 $X=107450 $Y=108560
X260 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=120980 106080 1 0 $X=120790 $Y=103120
X261 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=125120 122400 1 0 $X=124930 $Y=119440
X262 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=129720 95200 1 0 $X=129530 $Y=92240
X263 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=129720 155040 1 0 $X=129530 $Y=152080
X264 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=134780 51680 1 0 $X=134590 $Y=48720
X265 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=138460 89760 1 0 $X=138270 $Y=86800
X266 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=138920 68000 1 0 $X=138730 $Y=65040
X267 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=141680 62560 1 0 $X=141490 $Y=59600
X268 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=149960 100640 1 0 $X=149770 $Y=97680
X269 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=149960 122400 1 0 $X=149770 $Y=119440
X270 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4 $T=150420 29920 1 0 $X=150230 $Y=26960
X271 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 19040 0 0 $X=6710 $Y=18800
X272 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 116960 0 0 $X=6710 $Y=116720
X273 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 144160 1 0 $X=6710 $Y=141200
X274 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=6900 149600 1 0 $X=6710 $Y=146640
X275 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=11500 111520 1 0 $X=11310 $Y=108560
X276 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=16560 78880 1 0 $X=16370 $Y=75920
X277 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=17020 29920 1 0 $X=16830 $Y=26960
X278 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=17020 116960 0 0 $X=16830 $Y=116720
X279 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=20240 106080 1 0 $X=20050 $Y=103120
X280 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=22080 24480 1 0 $X=21890 $Y=21520
X281 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=22080 127840 1 0 $X=21890 $Y=124880
X282 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=31280 155040 0 0 $X=31090 $Y=154800
X283 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=31740 122400 1 0 $X=31550 $Y=119440
X284 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=34040 78880 0 0 $X=33850 $Y=78640
X285 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=39560 35360 0 0 $X=39370 $Y=35120
X286 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=39560 111520 0 0 $X=39370 $Y=111280
X287 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=44620 29920 1 0 $X=44430 $Y=26960
X288 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=45080 95200 1 0 $X=44890 $Y=92240
X289 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=45080 100640 1 0 $X=44890 $Y=97680
X290 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=48300 84320 1 0 $X=48110 $Y=81360
X291 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=51980 111520 1 0 $X=51790 $Y=108560
X292 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=52440 95200 1 0 $X=52250 $Y=92240
X293 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=53360 57120 1 0 $X=53170 $Y=54160
X294 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=55200 127840 1 0 $X=55010 $Y=124880
X295 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=62100 100640 0 0 $X=61910 $Y=100400
X296 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=65320 73440 1 0 $X=65130 $Y=70480
X297 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=66240 35360 0 0 $X=66050 $Y=35120
X298 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=73140 78880 1 0 $X=72950 $Y=75920
X299 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=73140 155040 1 0 $X=72950 $Y=152080
X300 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=78660 127840 1 0 $X=78470 $Y=124880
X301 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=78660 133280 1 0 $X=78470 $Y=130320
X302 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=78660 138720 1 0 $X=78470 $Y=135760
X303 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=81420 62560 1 0 $X=81230 $Y=59600
X304 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=83260 78880 1 0 $X=83070 $Y=75920
X305 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=84180 68000 1 0 $X=83990 $Y=65040
X306 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=85100 138720 1 0 $X=84910 $Y=135760
X307 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=86480 19040 1 0 $X=86290 $Y=16080
X308 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=86940 116960 1 0 $X=86750 $Y=114000
X309 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=90160 46240 1 0 $X=89970 $Y=43280
X310 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=90160 84320 0 0 $X=89970 $Y=84080
X311 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=92000 89760 0 0 $X=91810 $Y=89520
X312 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=96140 138720 1 0 $X=95950 $Y=135760
X313 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=96600 106080 1 0 $X=96410 $Y=103120
X314 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=97060 57120 1 0 $X=96870 $Y=54160
X315 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=97520 51680 0 0 $X=97330 $Y=51440
X316 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=100740 144160 1 0 $X=100550 $Y=141200
X317 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=103500 106080 0 0 $X=103310 $Y=105840
X318 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=104420 116960 1 0 $X=104230 $Y=114000
X319 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=107640 13600 1 0 $X=107450 $Y=10640
X320 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=108560 62560 0 0 $X=108370 $Y=62320
X321 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=109480 40800 1 0 $X=109290 $Y=37840
X322 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=109940 89760 1 0 $X=109750 $Y=86800
X323 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=110860 62560 1 0 $X=110670 $Y=59600
X324 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=119140 57120 1 0 $X=118950 $Y=54160
X325 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=120060 100640 1 0 $X=119870 $Y=97680
X326 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=129260 100640 1 0 $X=129070 $Y=97680
X327 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=132480 29920 1 0 $X=132290 $Y=26960
X328 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=132480 35360 1 0 $X=132290 $Y=32400
X329 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=132480 40800 1 0 $X=132290 $Y=37840
X330 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=132480 100640 1 0 $X=132290 $Y=97680
X331 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=134780 78880 1 0 $X=134590 $Y=75920
X332 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=136160 84320 1 0 $X=135970 $Y=81360
X333 VSS VDD VSS VDD sky130_fd_sc_hd__decap_6 $T=149040 111520 1 0 $X=148850 $Y=108560
X334 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=6900 78880 0 0 $X=6710 $Y=78640
X335 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=6900 133280 0 0 $X=6710 $Y=133040
X336 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=6900 138720 1 0 $X=6710 $Y=135760
X337 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=6900 155040 1 0 $X=6710 $Y=152080
X338 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=14260 24480 0 0 $X=14070 $Y=24240
X339 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=14720 155040 1 0 $X=14530 $Y=152080
X340 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=15180 68000 1 0 $X=14990 $Y=65040
X341 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=15180 144160 0 0 $X=14990 $Y=143920
X342 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=15640 144160 1 0 $X=15450 $Y=141200
X343 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=18400 73440 0 0 $X=18210 $Y=73200
X344 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=20240 13600 1 0 $X=20050 $Y=10640
X345 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=20240 19040 1 0 $X=20050 $Y=16080
X346 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=20240 73440 1 0 $X=20050 $Y=70480
X347 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=20240 149600 1 0 $X=20050 $Y=146640
X348 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=20240 155040 1 0 $X=20050 $Y=152080
X349 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=22080 35360 1 0 $X=21890 $Y=32400
X350 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=24380 122400 1 0 $X=24190 $Y=119440
X351 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=29440 106080 1 0 $X=29250 $Y=103120
X352 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43700 35360 1 0 $X=43510 $Y=32400
X353 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43700 106080 1 0 $X=43510 $Y=103120
X354 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=43700 111520 1 0 $X=43510 $Y=108560
X355 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=44160 133280 1 0 $X=43970 $Y=130320
X356 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=44620 68000 0 0 $X=44430 $Y=67760
X357 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=45080 62560 0 0 $X=44890 $Y=62320
X358 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=45540 78880 0 0 $X=45350 $Y=78640
X359 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=50140 89760 1 0 $X=49950 $Y=86800
X360 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=53820 78880 1 0 $X=53630 $Y=75920
X361 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=57500 57120 0 0 $X=57310 $Y=56880
X362 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=60720 116960 1 0 $X=60530 $Y=114000
X363 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=63020 46240 1 0 $X=62830 $Y=43280
X364 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=63020 111520 1 0 $X=62830 $Y=108560
X365 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=65320 100640 1 0 $X=65130 $Y=97680
X366 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=68080 29920 1 0 $X=67890 $Y=26960
X367 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=70840 138720 1 0 $X=70650 $Y=135760
X368 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=70840 144160 1 0 $X=70650 $Y=141200
X369 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=74060 138720 0 0 $X=73870 $Y=138480
X370 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=78200 68000 1 0 $X=78010 $Y=65040
X371 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=84640 51680 1 0 $X=84450 $Y=48720
X372 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=85560 62560 1 0 $X=85370 $Y=59600
X373 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=85560 106080 1 0 $X=85370 $Y=103120
X374 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=85560 111520 1 0 $X=85370 $Y=108560
X375 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=86480 149600 1 0 $X=86290 $Y=146640
X376 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=86940 122400 1 0 $X=86750 $Y=119440
X377 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=87400 144160 1 0 $X=87210 $Y=141200
X378 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=91080 57120 1 0 $X=90890 $Y=54160
X379 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=93380 111520 1 0 $X=93190 $Y=108560
X380 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=94760 89760 1 0 $X=94570 $Y=86800
X381 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=95220 13600 1 0 $X=95030 $Y=10640
X382 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=98900 84320 1 0 $X=98710 $Y=81360
X383 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=98900 116960 1 0 $X=98710 $Y=114000
X384 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=99820 40800 1 0 $X=99630 $Y=37840
X385 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=100280 95200 1 0 $X=100090 $Y=92240
X386 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=109480 73440 1 0 $X=109290 $Y=70480
X387 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=113160 35360 1 0 $X=112970 $Y=32400
X388 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=113620 40800 1 0 $X=113430 $Y=37840
X389 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=113620 122400 1 0 $X=113430 $Y=119440
X390 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=113620 127840 1 0 $X=113430 $Y=124880
X391 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=116380 144160 1 0 $X=116190 $Y=141200
X392 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=119600 73440 1 0 $X=119410 $Y=70480
X393 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=122360 127840 0 0 $X=122170 $Y=127600
X394 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=123740 144160 1 0 $X=123550 $Y=141200
X395 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=126960 19040 1 0 $X=126770 $Y=16080
X396 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=128340 51680 1 0 $X=128150 $Y=48720
X397 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=132480 111520 1 0 $X=132290 $Y=108560
X398 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=134320 155040 1 0 $X=134130 $Y=152080
X399 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=142600 35360 1 0 $X=142410 $Y=32400
X400 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=147660 35360 1 0 $X=147470 $Y=32400
X401 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=147660 68000 1 0 $X=147470 $Y=65040
X402 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8 $T=148580 127840 1 0 $X=148390 $Y=124880
X453 VSS VDD ICV_4 $T=47840 24480 1 0 $X=47650 $Y=21520
X454 VSS VDD ICV_4 $T=61640 13600 0 0 $X=61450 $Y=13360
X455 VSS VDD ICV_4 $T=61640 57120 0 0 $X=61450 $Y=56880
X456 VSS VDD ICV_4 $T=75900 122400 1 0 $X=75710 $Y=119440
X457 VSS VDD ICV_4 $T=89700 57120 0 0 $X=89510 $Y=56880
X458 VSS VDD ICV_4 $T=91080 155040 0 0 $X=90890 $Y=154800
X459 VSS VDD ICV_4 $T=103960 24480 1 0 $X=103770 $Y=21520
X460 VSS VDD ICV_4 $T=103960 138720 1 0 $X=103770 $Y=135760
X461 VSS VDD ICV_4 $T=132020 46240 1 0 $X=131830 $Y=43280
X462 VSS VDD ICV_4 $T=148120 13600 1 0 $X=147930 $Y=10640
X463 VSS VDD ICV_4 $T=148120 155040 0 0 $X=147930 $Y=154800
X464 VSS VDD ICV_5 $T=148120 78880 1 0 $X=147930 $Y=75920
X465 VSS VDD ICV_6 $T=15180 138720 0 0 $X=14990 $Y=138480
X466 VSS VDD ICV_6 $T=22540 111520 1 0 $X=22350 $Y=108560
X467 VSS VDD ICV_6 $T=34960 133280 1 0 $X=34770 $Y=130320
X468 VSS VDD ICV_6 $T=70840 116960 1 0 $X=70650 $Y=114000
X469 VSS VDD ICV_6 $T=124200 144160 0 0 $X=124010 $Y=143920
X470 VSS VDD ICV_6 $T=126960 40800 0 0 $X=126770 $Y=40560
X471 VSS VDD ICV_6 $T=140760 106080 0 0 $X=140570 $Y=105840
X472 VSS VDD ICV_6 $T=140760 149600 0 0 $X=140570 $Y=149360
X473 VSS VDD ICV_6 $T=147200 46240 1 0 $X=147010 $Y=43280
X474 VSS VDD ICV_6 $T=147200 138720 1 0 $X=147010 $Y=135760
X475 VSS VDD ICV_6 $T=147200 144160 1 0 $X=147010 $Y=141200
X476 VSS VDD ICV_6 $T=147200 149600 1 0 $X=147010 $Y=146640
X477 VSS RESET sky130_fd_sc_hd__diode_2 $T=11500 35360 0 0 $X=11310 $Y=35120
X478 VSS 100 sky130_fd_sc_hd__diode_2 $T=12420 95200 0 0 $X=12230 $Y=94960
X479 VSS 155 sky130_fd_sc_hd__diode_2 $T=23460 106080 1 0 $X=23270 $Y=103120
X480 VSS 133 sky130_fd_sc_hd__diode_2 $T=23920 68000 0 0 $X=23730 $Y=67760
X481 VSS 222 sky130_fd_sc_hd__diode_2 $T=37720 84320 0 0 $X=37530 $Y=84080
X482 VSS 56 sky130_fd_sc_hd__diode_2 $T=38180 46240 1 0 $X=37990 $Y=43280
X483 VSS COUNT<0> sky130_fd_sc_hd__diode_2 $T=42320 89760 0 0 $X=42130 $Y=89520
X484 VSS SAMPLE_COUNT<2> sky130_fd_sc_hd__diode_2 $T=44620 51680 0 0 $X=44430 $Y=51440
X485 VSS 242 sky130_fd_sc_hd__diode_2 $T=45540 111520 0 0 $X=45350 $Y=111280
X486 VSS 118 sky130_fd_sc_hd__diode_2 $T=51520 122400 1 0 $X=51330 $Y=119440
X487 VSS 281 sky130_fd_sc_hd__diode_2 $T=51520 127840 0 0 $X=51330 $Y=127600
X488 VSS 217 sky130_fd_sc_hd__diode_2 $T=52900 116960 1 0 $X=52710 $Y=114000
X489 VSS 306 sky130_fd_sc_hd__diode_2 $T=55200 111520 1 0 $X=55010 $Y=108560
X490 VSS PAR_IN1<7> sky130_fd_sc_hd__diode_2 $T=66700 78880 0 0 $X=66510 $Y=78640
X491 VSS 385 sky130_fd_sc_hd__diode_2 $T=67620 95200 0 0 $X=67430 $Y=94960
X492 VSS 396 sky130_fd_sc_hd__diode_2 $T=68080 138720 0 0 $X=67890 $Y=138480
X493 VSS 383 sky130_fd_sc_hd__diode_2 $T=80040 127840 0 0 $X=79850 $Y=127600
X494 VSS 272 sky130_fd_sc_hd__diode_2 $T=81420 19040 1 0 $X=81230 $Y=16080
X495 VSS 497 sky130_fd_sc_hd__diode_2 $T=87400 68000 1 0 $X=87210 $Y=65040
X496 VSS 392 sky130_fd_sc_hd__diode_2 $T=97520 29920 0 0 $X=97330 $Y=29680
X497 VSS 567 sky130_fd_sc_hd__diode_2 $T=97520 106080 0 0 $X=97330 $Y=105840
X498 VSS 650 sky130_fd_sc_hd__diode_2 $T=113620 73440 1 0 $X=113430 $Y=70480
X499 VSS 290 sky130_fd_sc_hd__diode_2 $T=122360 51680 1 0 $X=122170 $Y=48720
X500 VSS 56 75 ICV_7 $T=7820 35360 0 0 $X=7630 $Y=35120
X501 VSS RESET READY ICV_7 $T=7820 57120 0 0 $X=7630 $Y=56880
X502 VSS PAR_IN7<13> 77 ICV_7 $T=7820 84320 0 0 $X=7630 $Y=84080
X503 VSS PAR_IN7<29> 77 ICV_7 $T=7820 116960 1 0 $X=7630 $Y=114000
X504 VSS PAR_IN6<29> 59 ICV_7 $T=8280 106080 0 0 $X=8090 $Y=105840
X505 VSS 49 RESET ICV_7 $T=9660 19040 0 0 $X=9470 $Y=18800
X506 VSS PAR_IN4<4> 80 ICV_7 $T=10580 133280 0 0 $X=10390 $Y=133040
X507 VSS PAR_IN6<25> 103 ICV_7 $T=12420 138720 0 0 $X=12230 $Y=138480
X508 VSS 7 4 ICV_7 $T=12880 51680 0 0 $X=12690 $Y=51440
X509 VSS 100 14 ICV_7 $T=14260 89760 1 0 $X=14070 $Y=86800
X510 VSS 107 109 ICV_7 $T=14260 95200 1 0 $X=14070 $Y=92240
X511 VSS 115 56 ICV_7 $T=16100 46240 1 0 $X=15910 $Y=43280
X512 VSS 116 97 ICV_7 $T=16560 84320 0 0 $X=16370 $Y=84080
X513 VSS 83 COUNT<5> ICV_7 $T=18400 24480 0 0 $X=18210 $Y=24240
X514 VSS COMPLETE 135 ICV_7 $T=19780 78880 0 0 $X=19590 $Y=78640
X515 VSS 89 PAR_IN8<21> ICV_7 $T=20240 13600 0 0 $X=20050 $Y=13360
X516 VSS 129 140 ICV_7 $T=20240 138720 0 0 $X=20050 $Y=138480
X517 VSS 136 154 ICV_7 $T=21620 100640 1 0 $X=21430 $Y=97680
X518 VSS READY COMPLETE ICV_7 $T=23000 57120 0 0 $X=22810 $Y=56880
X519 VSS 69 12 ICV_7 $T=24380 57120 1 0 $X=24190 $Y=54160
X520 VSS PAR_IN8<13> 146 ICV_7 $T=26680 73440 0 0 $X=26490 $Y=73200
X521 VSS 146 COUNT<5> ICV_7 $T=28060 62560 0 0 $X=27870 $Y=62320
X522 VSS PAR_IN5<8> 102 ICV_7 $T=29900 138720 0 0 $X=29710 $Y=138480
X523 VSS 12 211 ICV_7 $T=34500 46240 1 0 $X=34310 $Y=43280
X524 VSS 6 205 ICV_7 $T=34960 24480 0 0 $X=34770 $Y=24240
X525 VSS 181 PAR_IN4<20> ICV_7 $T=36340 13600 0 0 $X=36150 $Y=13360
X526 VSS 188 238 ICV_7 $T=40020 138720 1 0 $X=39830 $Y=135760
X527 VSS 239 215 ICV_7 $T=42780 46240 0 0 $X=42590 $Y=46000
X528 VSS 184 SAMPLE_COUNT<2> ICV_7 $T=43240 40800 0 0 $X=43050 $Y=40560
X529 VSS 143 184 ICV_7 $T=45080 57120 0 0 $X=44890 $Y=56880
X530 VSS 18 COUNT<2> ICV_7 $T=45080 95200 0 0 $X=44890 $Y=94960
X531 VSS 252 14 ICV_7 $T=46000 106080 0 0 $X=45810 $Y=105840
X532 VSS 256 261 ICV_7 $T=46460 73440 0 0 $X=46270 $Y=73200
X533 VSS 273 PAR_IN3<5> ICV_7 $T=49680 78880 0 0 $X=49490 $Y=78640
X534 VSS 265 240 ICV_7 $T=51520 40800 1 0 $X=51330 $Y=37840
X535 VSS 279 291 ICV_7 $T=51520 100640 1 0 $X=51330 $Y=97680
X536 VSS PAR_IN1<24> 281 ICV_7 $T=53820 116960 0 0 $X=53630 $Y=116720
X537 VSS 207 112 ICV_7 $T=54740 29920 0 0 $X=54550 $Y=29680
X538 VSS SAMPLE_COUNT<2> 184 ICV_7 $T=56120 51680 0 0 $X=55930 $Y=51440
X539 VSS 18 18 ICV_7 $T=56120 89760 0 0 $X=55930 $Y=89520
X540 VSS PAR_IN7<6> 286 ICV_7 $T=57500 73440 0 0 $X=57310 $Y=73200
X541 VSS PAR_IN1<9> 262 ICV_7 $T=57500 127840 0 0 $X=57310 $Y=127600
X542 VSS 323 203 ICV_7 $T=57960 127840 1 0 $X=57770 $Y=124880
X543 VSS 211 268 ICV_7 $T=58880 40800 1 0 $X=58690 $Y=37840
X544 VSS PAR_IN3<7> 289 ICV_7 $T=63020 19040 0 0 $X=62830 $Y=18800
X545 VSS PAR_IN2<9> PAR_IN3<24> ICV_7 $T=63020 133280 0 0 $X=62830 $Y=133040
X546 VSS 229 262 ICV_7 $T=63940 62560 0 0 $X=63750 $Y=62320
X547 VSS COUNT<3> PAR_IN2<14> ICV_7 $T=64400 111520 0 0 $X=64210 $Y=111280
X548 VSS 127 PAR_IN5<2> ICV_7 $T=64860 40800 1 0 $X=64670 $Y=37840
X549 VSS 365 COUNT<2> ICV_7 $T=65320 100640 0 0 $X=65130 $Y=100400
X550 VSS 351 383 ICV_7 $T=65320 144160 1 0 $X=65130 $Y=141200
X551 VSS 229 387 ICV_7 $T=65780 133280 1 0 $X=65590 $Y=130320
X552 VSS 408 118 ICV_7 $T=71300 68000 0 0 $X=71110 $Y=67760
X553 VSS 411 14 ICV_7 $T=71300 84320 0 0 $X=71110 $Y=84080
X554 VSS 377 418 ICV_7 $T=71760 29920 1 0 $X=71570 $Y=26960
X555 VSS 413 PAR_IN1<31> ICV_7 $T=72220 13600 0 0 $X=72030 $Y=13360
X556 VSS 414 421 ICV_7 $T=72220 35360 1 0 $X=72030 $Y=32400
X557 VSS 416 373 ICV_7 $T=72680 57120 0 0 $X=72490 $Y=56880
X558 VSS 430 448 ICV_7 $T=76360 95200 0 0 $X=76170 $Y=94960
X559 VSS 206 341 ICV_7 $T=76360 127840 0 0 $X=76170 $Y=127600
X560 VSS 341 395 ICV_7 $T=77740 122400 0 0 $X=77550 $Y=122160
X561 VSS 203 451 ICV_7 $T=77740 138720 0 0 $X=77550 $Y=138480
X562 VSS 450 457 ICV_7 $T=78200 111520 0 0 $X=78010 $Y=111280
X563 VSS 348 465 ICV_7 $T=79580 73440 1 0 $X=79390 $Y=70480
X564 VSS 118 483 ICV_7 $T=81880 84320 0 0 $X=81690 $Y=84080
X565 VSS 468 77 ICV_7 $T=83720 24480 1 0 $X=83530 $Y=21520
X566 VSS PAR_IN1<22> 303 ICV_7 $T=83720 116960 0 0 $X=83530 $Y=116720
X567 VSS 487 135 ICV_7 $T=86020 73440 0 0 $X=85830 $Y=73200
X568 VSS 493 PAR_IN6<20> ICV_7 $T=86020 100640 0 0 $X=85830 $Y=100400
X569 VSS 495 505 ICV_7 $T=86480 78880 1 0 $X=86290 $Y=75920
X570 VSS 507 478 ICV_7 $T=88320 133280 1 0 $X=88130 $Y=130320
X571 VSS 508 281 ICV_7 $T=88320 138720 1 0 $X=88130 $Y=135760
X572 VSS PAR_IN2<29> 336 ICV_7 $T=93380 40800 0 0 $X=93190 $Y=40560
X573 VSS PAR_IN3<6> 228 ICV_7 $T=94760 89760 0 0 $X=94570 $Y=89520
X574 VSS 288 547 ICV_7 $T=95220 78880 1 0 $X=95030 $Y=75920
X575 VSS PAR_IN1<17> PAR_IN1<27> ICV_7 $T=96140 13600 0 0 $X=95950 $Y=13360
X576 VSS PAR_IN8<1> 524 ICV_7 $T=97060 116960 0 0 $X=96870 $Y=116720
X577 VSS PAR_IN7<5> 575 ICV_7 $T=100280 149600 1 0 $X=100090 $Y=146640
X578 VSS PAR_IN1<3> PAR_IN6<28> ICV_7 $T=103960 13600 0 0 $X=103770 $Y=13360
X579 VSS PAR_IN5<19> 563 ICV_7 $T=104420 40800 0 0 $X=104230 $Y=40560
X580 VSS PAR_IN3<3> 91 ICV_7 $T=106260 57120 0 0 $X=106070 $Y=56880
X581 VSS 610 374 ICV_7 $T=106260 95200 0 0 $X=106070 $Y=94960
X582 VSS 556 622 ICV_7 $T=106260 106080 0 0 $X=106070 $Y=105840
X583 VSS 558 606 ICV_7 $T=108100 138720 1 0 $X=107910 $Y=135760
X584 VSS 629 164 ICV_7 $T=109480 19040 1 0 $X=109290 $Y=16080
X585 VSS 626 PAR_IN8<11> ICV_7 $T=111780 62560 0 0 $X=111590 $Y=62320
X586 VSS PAR_IN3<10> PAR_IN5<10> ICV_7 $T=111780 89760 0 0 $X=111590 $Y=89520
X587 VSS PAR_IN6<3> 643 ICV_7 $T=113160 13600 1 0 $X=112970 $Y=10640
X588 VSS 653 PAR_IN4<19> ICV_7 $T=114080 78880 0 0 $X=113890 $Y=78640
X589 VSS 668 672 ICV_7 $T=116380 116960 1 0 $X=116190 $Y=114000
X590 VSS 604 PAR_IN3<26> ICV_7 $T=119140 100640 0 0 $X=118950 $Y=100400
X591 VSS PAR_IN4<9> 602 ICV_7 $T=121440 144160 0 0 $X=121250 $Y=143920
X592 VSS 674 706 ICV_7 $T=124200 40800 0 0 $X=124010 $Y=40560
X593 VSS 709 729 ICV_7 $T=126500 57120 1 0 $X=126310 $Y=54160
X594 VSS 620 546 ICV_7 $T=127880 19040 0 0 $X=127690 $Y=18800
X595 VSS 726 727 ICV_7 $T=127880 111520 1 0 $X=127690 $Y=108560
X596 VSS 698 707 ICV_7 $T=127880 116960 1 0 $X=127690 $Y=114000
X597 VSS 731 510 ICV_7 $T=128340 68000 1 0 $X=128150 $Y=65040
X598 VSS PAR_IN5<16> PAR_IN6<27> ICV_7 $T=132480 13600 0 0 $X=132290 $Y=13360
X599 VSS PAR_IN8<18> 329 ICV_7 $T=132940 51680 0 0 $X=132750 $Y=51440
X600 VSS PAR_IN2<18> 654 ICV_7 $T=133860 62560 0 0 $X=133670 $Y=62320
X601 VSS PAR_IN5<30> 289 ICV_7 $T=135700 40800 1 0 $X=135510 $Y=37840
X602 VSS 767 780 ICV_7 $T=142140 29920 0 0 $X=141950 $Y=29680
X603 VSS 620 776 ICV_7 $T=142140 40800 0 0 $X=141950 $Y=40560
X604 VSS VDD 65 82 ICV_8 $T=8280 51680 0 0 $X=8090 $Y=51440
X605 VSS VDD 89 PAR_IN5<29> ICV_8 $T=11040 78880 0 0 $X=10850 $Y=78640
X606 VSS VDD 116 152 ICV_8 $T=21160 78880 1 0 $X=20970 $Y=75920
X607 VSS VDD 143 6 ICV_8 $T=22540 40800 1 0 $X=22350 $Y=37840
X608 VSS VDD PAR_IN1<12> 186 ICV_8 $T=28520 116960 0 0 $X=28330 $Y=116720
X609 VSS VDD 178 156 ICV_8 $T=28520 133280 0 0 $X=28330 $Y=133040
X610 VSS VDD 190 165 ICV_8 $T=34040 19040 1 0 $X=33850 $Y=16080
X611 VSS VDD 82 192 ICV_8 $T=34960 40800 0 0 $X=34770 $Y=40560
X612 VSS VDD 206 195 ICV_8 $T=34960 122400 1 0 $X=34770 $Y=119440
X613 VSS VDD PAR_IN1<8> 186 ICV_8 $T=35880 133280 0 0 $X=35690 $Y=133040
X614 VSS VDD 258 PAR_IN2<12> ICV_8 $T=46460 138720 0 0 $X=46270 $Y=138480
X615 VSS VDD PAR_IN6<4> 103 ICV_8 $T=49220 149600 1 0 $X=49030 $Y=146640
X616 VSS VDD 215 211 ICV_8 $T=51520 51680 0 0 $X=51330 $Y=51440
X617 VSS VDD PAR_IN1<2> 303 ICV_8 $T=56580 62560 0 0 $X=56390 $Y=62320
X618 VSS VDD 258 PAR_IN2<16> ICV_8 $T=56580 100640 0 0 $X=56390 $Y=100400
X619 VSS VDD 262 317 ICV_8 $T=61180 68000 1 0 $X=60990 $Y=65040
X620 VSS VDD 71 348 ICV_8 $T=70840 40800 1 0 $X=70650 $Y=37840
X621 VSS VDD 432 390 ICV_8 $T=77280 29920 1 0 $X=77090 $Y=26960
X622 VSS VDD 413 472 ICV_8 $T=83720 133280 1 0 $X=83530 $Y=130320
X623 VSS VDD PAR_IN1<15> 281 ICV_8 $T=84640 133280 0 0 $X=84450 $Y=133040
X624 VSS VDD 447 469 ICV_8 $T=85100 89760 0 0 $X=84910 $Y=89520
X625 VSS VDD 431 PAR_IN4<5> ICV_8 $T=89700 19040 1 0 $X=89510 $Y=16080
X626 VSS VDD 202 527 ICV_8 $T=90160 73440 1 0 $X=89970 $Y=70480
X627 VSS VDD PAR_IN4<24> 80 ICV_8 $T=91080 144160 0 0 $X=90890 $Y=143920
X628 VSS VDD 530 538 ICV_8 $T=92000 133280 1 0 $X=91810 $Y=130320
X629 VSS VDD PAR_IN4<15> 59 ICV_8 $T=101200 95200 0 0 $X=101010 $Y=94960
X630 VSS VDD 432 630 ICV_8 $T=108560 24480 1 0 $X=108370 $Y=21520
X631 VSS VDD PAR_IN3<30> 457 ICV_8 $T=119140 40800 0 0 $X=118950 $Y=40560
X632 VSS VDD 282 77 ICV_8 $T=123280 68000 1 0 $X=123090 $Y=65040
X633 VSS VDD PAR_IN6<31> 643 ICV_8 $T=123740 13600 0 0 $X=123550 $Y=13360
X634 VSS VDD 672 747 ICV_8 $T=133860 127840 0 0 $X=133670 $Y=127600
X635 VSS VDD PAR_IN4<30> PAR_IN2<27> ICV_8 $T=141220 46240 0 0 $X=141030 $Y=46000
X636 VSS VDD PAR_IN2<23> 272 ICV_8 $T=147200 73440 0 0 $X=147010 $Y=73200
X637 VSS VDD 145 795 ICV_8 $T=147200 89760 0 0 $X=147010 $Y=89520
X638 VSS VDD 387 788 ICV_8 $T=147200 133280 0 0 $X=147010 $Y=133040
X639 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 13600 0 0 $X=6710 $Y=13360
X640 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 19040 1 0 $X=6710 $Y=16080
X641 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 24480 1 0 $X=6710 $Y=21520
X642 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 84320 1 0 $X=6710 $Y=81360
X643 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 95200 0 0 $X=6710 $Y=94960
X644 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=6900 138720 0 0 $X=6710 $Y=138480
X645 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=14260 68000 0 0 $X=14070 $Y=67760
X646 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=24840 127840 0 0 $X=24650 $Y=127600
X647 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=27140 111520 0 0 $X=26950 $Y=111280
X648 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=37260 149600 1 0 $X=37070 $Y=146640
X649 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=37720 100640 0 0 $X=37530 $Y=100400
X650 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=38180 111520 1 0 $X=37990 $Y=108560
X651 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=38180 127840 1 0 $X=37990 $Y=124880
X652 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=39560 106080 0 0 $X=39370 $Y=105840
X653 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=40480 62560 1 0 $X=40290 $Y=59600
X654 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=40480 84320 1 0 $X=40290 $Y=81360
X655 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=47840 144160 0 0 $X=47650 $Y=143920
X656 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=50140 84320 0 0 $X=49950 $Y=84080
X657 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=53820 35360 0 0 $X=53630 $Y=35120
X658 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=56580 122400 1 0 $X=56390 $Y=119440
X659 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=57960 62560 1 0 $X=57770 $Y=59600
X660 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=60260 57120 1 0 $X=60070 $Y=54160
X661 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=60720 155040 1 0 $X=60530 $Y=152080
X662 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=63480 95200 1 0 $X=63290 $Y=92240
X663 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=64400 122400 1 0 $X=64210 $Y=119440
X664 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69460 51680 1 0 $X=69270 $Y=48720
X665 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69460 57120 1 0 $X=69270 $Y=54160
X666 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69920 24480 1 0 $X=69730 $Y=21520
X667 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=69920 89760 1 0 $X=69730 $Y=86800
X668 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=70380 68000 1 0 $X=70190 $Y=65040
X669 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=80040 106080 1 0 $X=79850 $Y=103120
X670 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=81880 144160 1 0 $X=81690 $Y=141200
X671 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=83720 84320 1 0 $X=83530 $Y=81360
X672 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=84640 13600 1 0 $X=84450 $Y=10640
X673 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=95220 68000 1 0 $X=95030 $Y=65040
X674 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=96600 73440 1 0 $X=96410 $Y=70480
X675 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=108100 122400 1 0 $X=107910 $Y=119440
X676 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=108560 155040 1 0 $X=108370 $Y=152080
X677 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=110860 84320 1 0 $X=110670 $Y=81360
X678 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=112700 133280 1 0 $X=112510 $Y=130320
X679 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=113160 138720 1 0 $X=112970 $Y=135760
X680 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=121900 35360 0 0 $X=121710 $Y=35120
X681 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=122360 19040 0 0 $X=122170 $Y=18800
X682 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=122820 40800 1 0 $X=122630 $Y=37840
X683 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=136160 62560 1 0 $X=135970 $Y=59600
X684 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=141680 46240 1 0 $X=141490 $Y=43280
X685 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=141680 144160 1 0 $X=141490 $Y=141200
X686 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=145360 57120 1 0 $X=145170 $Y=54160
X687 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=145820 40800 1 0 $X=145630 $Y=37840
X688 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=145820 95200 1 0 $X=145630 $Y=92240
X689 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146280 62560 0 0 $X=146090 $Y=62320
X690 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146280 68000 0 0 $X=146090 $Y=67760
X691 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146280 78880 0 0 $X=146090 $Y=78640
X692 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146280 133280 1 0 $X=146090 $Y=130320
X693 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146740 73440 1 0 $X=146550 $Y=70480
X694 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12 $T=146740 84320 1 0 $X=146550 $Y=81360
X695 VSS VDD SAMPLE_COUNT<2> VDD 56 VSS sky130_fd_sc_hd__buf_1 $T=7820 46240 1 0 $X=7630 $Y=43280
X696 VSS VDD 103 VDD 59 VSS sky130_fd_sc_hd__buf_1 $T=15180 122400 0 0 $X=14990 $Y=122160
X697 VSS VDD 113 VDD 82 VSS sky130_fd_sc_hd__buf_1 $T=22080 62560 0 0 $X=21890 $Y=62320
X698 VSS VDD COMPLETE VDD 6 VSS sky130_fd_sc_hd__buf_1 $T=26680 57120 0 0 $X=26490 $Y=56880
X699 VSS VDD 166 VDD 133 VSS sky130_fd_sc_hd__buf_1 $T=26680 78880 0 0 $X=26490 $Y=78640
X700 VSS VDD 203 VDD 135 VSS sky130_fd_sc_hd__buf_1 $T=35880 116960 0 0 $X=35690 $Y=116720
X701 VSS VDD 215 VDD 69 VSS sky130_fd_sc_hd__buf_1 $T=37720 57120 0 0 $X=37530 $Y=56880
X702 VSS VDD 239 VDD 215 VSS sky130_fd_sc_hd__buf_1 $T=42780 51680 1 0 $X=42590 $Y=48720
X703 VSS VDD 18 VDD 14 VSS sky130_fd_sc_hd__buf_1 $T=53820 89760 0 0 $X=53630 $Y=89520
X704 VSS VDD 262 VDD 227 VSS sky130_fd_sc_hd__buf_1 $T=53820 133280 0 0 $X=53630 $Y=133040
X705 VSS VDD SAMPLE_COUNT<0> VDD 184 VSS sky130_fd_sc_hd__buf_1 $T=54740 40800 0 0 $X=54550 $Y=40560
X706 VSS VDD 258 VDD 272 VSS sky130_fd_sc_hd__buf_1 $T=54740 73440 1 0 $X=54550 $Y=70480
X707 VSS VDD 262 VDD 203 VSS sky130_fd_sc_hd__buf_1 $T=55660 133280 1 0 $X=55470 $Y=130320
X708 VSS VDD 319 VDD 202 VSS sky130_fd_sc_hd__buf_1 $T=63020 89760 0 0 $X=62830 $Y=89520
X709 VSS VDD COUNT<3> VDD 319 VSS sky130_fd_sc_hd__buf_1 $T=64400 116960 1 0 $X=64210 $Y=114000
X710 VSS VDD 301 VDD 228 VSS sky130_fd_sc_hd__buf_1 $T=66240 57120 0 0 $X=66050 $Y=56880
X711 VSS VDD COUNT<4> VDD 341 VSS sky130_fd_sc_hd__buf_1 $T=69460 127840 1 0 $X=69270 $Y=124880
X712 VSS VDD 348 VDD 207 VSS sky130_fd_sc_hd__buf_1 $T=72680 40800 0 0 $X=72490 $Y=40560
X713 VSS VDD 348 VDD 102 VSS sky130_fd_sc_hd__buf_1 $T=75900 62560 0 0 $X=75710 $Y=62320
X714 VSS VDD 373 VDD 348 VSS sky130_fd_sc_hd__buf_1 $T=76360 57120 0 0 $X=76170 $Y=56880
X715 VSS VDD 281 VDD 401 VSS sky130_fd_sc_hd__buf_1 $T=76360 116960 0 0 $X=76170 $Y=116720
X716 VSS VDD 383 VDD 281 VSS sky130_fd_sc_hd__buf_1 $T=77280 138720 1 0 $X=77090 $Y=135760
X717 VSS VDD 383 VDD 413 VSS sky130_fd_sc_hd__buf_1 $T=81420 133280 1 0 $X=81230 $Y=130320
X718 VSS VDD 395 VDD 336 VSS sky130_fd_sc_hd__buf_1 $T=81880 127840 1 0 $X=81690 $Y=124880
X719 VSS VDD 329 VDD 373 VSS sky130_fd_sc_hd__buf_1 $T=84180 62560 1 0 $X=83990 $Y=59600
X720 VSS VDD 396 VDD 469 VSS sky130_fd_sc_hd__buf_1 $T=85560 46240 1 0 $X=85370 $Y=43280
X721 VSS VDD 228 VDD 91 VSS sky130_fd_sc_hd__buf_1 $T=95220 73440 1 0 $X=95030 $Y=70480
X722 VSS VDD 80 VDD 431 VSS sky130_fd_sc_hd__buf_1 $T=98440 127840 0 0 $X=98250 $Y=127600
X723 VSS VDD 556 VDD 81 VSS sky130_fd_sc_hd__buf_1 $T=101660 100640 0 0 $X=101470 $Y=100400
X724 VSS VDD 556 VDD 493 VSS sky130_fd_sc_hd__buf_1 $T=105340 106080 1 0 $X=105150 $Y=103120
X725 VSS VDD 602 VDD 80 VSS sky130_fd_sc_hd__buf_1 $T=105800 144160 1 0 $X=105610 $Y=141200
X726 VSS VDD 556 VDD 304 VSS sky130_fd_sc_hd__buf_1 $T=106260 111520 1 0 $X=106070 $Y=108560
X727 VSS VDD 282 VDD 395 VSS sky130_fd_sc_hd__buf_1 $T=107640 78880 0 0 $X=107450 $Y=78640
X728 VSS VDD 264 VDD 546 VSS sky130_fd_sc_hd__buf_1 $T=109480 35360 1 0 $X=109290 $Y=32400
X729 VSS VDD 374 VDD 556 VSS sky130_fd_sc_hd__buf_1 $T=109480 100640 1 0 $X=109290 $Y=97680
X730 VSS VDD 625 VDD 103 VSS sky130_fd_sc_hd__buf_1 $T=111780 138720 1 0 $X=111590 $Y=135760
X731 VSS VDD 264 VDD 625 VSS sky130_fd_sc_hd__buf_1 $T=112240 40800 1 0 $X=112050 $Y=37840
X732 VSS VDD 271 VDD 604 VSS sky130_fd_sc_hd__buf_1 $T=113620 62560 1 0 $X=113430 $Y=59600
X733 VSS VDD 558 VDD 164 VSS sky130_fd_sc_hd__buf_1 $T=115000 144160 1 0 $X=114810 $Y=141200
X734 VSS VDD 282 VDD 654 VSS sky130_fd_sc_hd__buf_1 $T=123280 73440 1 0 $X=123090 $Y=70480
X735 VSS VDD 654 VDD 290 VSS sky130_fd_sc_hd__buf_1 $T=127880 78880 0 0 $X=127690 $Y=78640
X736 VSS VDD 672 VDD 437 VSS sky130_fd_sc_hd__buf_1 $T=131560 127840 0 0 $X=131370 $Y=127600
X737 VSS VDD 677 VDD 77 VSS sky130_fd_sc_hd__buf_1 $T=132020 106080 0 0 $X=131830 $Y=105840
X738 VSS VDD 560 VDD 653 VSS sky130_fd_sc_hd__buf_1 $T=134320 106080 1 0 $X=134130 $Y=103120
X739 VSS VDD 285 VDD 617 VSS sky130_fd_sc_hd__buf_1 $T=134780 62560 1 0 $X=134590 $Y=59600
X740 VSS VDD 546 VDD 643 VSS sky130_fd_sc_hd__buf_1 $T=135700 24480 0 0 $X=135510 $Y=24240
X741 VSS VDD 140 VDD 89 VSS sky130_fd_sc_hd__buf_1 $T=137080 89760 1 0 $X=136890 $Y=86800
X742 VSS VDD 207 VDD 145 VSS sky130_fd_sc_hd__buf_1 $T=146280 35360 1 0 $X=146090 $Y=32400
X743 VSS VDD ICV_9 $T=33580 35360 0 0 $X=33390 $Y=35120
X744 VSS VDD ICV_9 $T=33580 106080 0 0 $X=33390 $Y=105840
X745 VSS VDD ICV_9 $T=33580 111520 0 0 $X=33390 $Y=111280
X746 VSS VDD ICV_9 $T=34040 13600 1 0 $X=33850 $Y=10640
X747 VSS VDD ICV_9 $T=47840 133280 1 0 $X=47650 $Y=130320
X748 VSS VDD ICV_9 $T=48300 13600 1 0 $X=48110 $Y=10640
X749 VSS VDD ICV_9 $T=61640 95200 0 0 $X=61450 $Y=94960
X750 VSS VDD ICV_9 $T=75900 116960 1 0 $X=75710 $Y=114000
X751 VSS VDD ICV_9 $T=103960 89760 1 0 $X=103770 $Y=86800
X752 VSS VDD ICV_9 $T=117760 62560 0 0 $X=117570 $Y=62320
X753 VSS VDD ICV_9 $T=132020 133280 1 0 $X=131830 $Y=130320
X754 VSS VDD ICV_9 $T=145820 24480 0 0 $X=145630 $Y=24240
X755 VSS VDD ICV_9 $T=145820 35360 0 0 $X=145630 $Y=35120
X756 VSS VDD ICV_9 $T=145820 40800 0 0 $X=145630 $Y=40560
X757 VSS VDD ICV_9 $T=145820 95200 0 0 $X=145630 $Y=94960
X758 VSS VDD ICV_9 $T=145820 100640 0 0 $X=145630 $Y=100400
X759 VSS VDD ICV_9 $T=145820 106080 0 0 $X=145630 $Y=105840
X760 VSS VDD ICV_9 $T=145820 111520 0 0 $X=145630 $Y=111280
X761 VSS VDD ICV_9 $T=145820 116960 0 0 $X=145630 $Y=116720
X762 VSS VDD ICV_9 $T=145820 122400 0 0 $X=145630 $Y=122160
X763 VSS VDD ICV_9 $T=145820 127840 0 0 $X=145630 $Y=127600
X764 VSS VDD ICV_9 $T=145820 138720 0 0 $X=145630 $Y=138480
X765 VSS VDD ICV_9 $T=145820 149600 0 0 $X=145630 $Y=149360
X766 VSS 97 ICV_10 $T=19780 24480 1 0 $X=19590 $Y=21520
X767 VSS 76 ICV_10 $T=19780 35360 1 0 $X=19590 $Y=32400
X768 VSS 127 ICV_10 $T=19780 127840 1 0 $X=19590 $Y=124880
X769 VSS 239 ICV_10 $T=47840 46240 1 0 $X=47650 $Y=43280
X770 VSS 130 ICV_10 $T=47840 51680 1 0 $X=47650 $Y=48720
X771 VSS 34 ICV_10 $T=47840 89760 1 0 $X=47650 $Y=86800
X772 VSS 409 ICV_10 $T=75900 68000 1 0 $X=75710 $Y=65040
X773 VSS PAR_IN3<14> ICV_10 $T=89700 46240 0 0 $X=89510 $Y=46000
X774 VSS 135 ICV_10 $T=89700 78880 0 0 $X=89510 $Y=78640
X775 VSS 492 ICV_10 $T=89700 89760 0 0 $X=89510 $Y=89520
X776 VSS 556 ICV_10 $T=103960 100640 1 0 $X=103770 $Y=97680
X777 VSS 546 ICV_10 $T=105340 13600 1 0 $X=105150 $Y=10640
X778 VSS PAR_IN7<1> ICV_10 $T=117760 116960 0 0 $X=117570 $Y=116720
X779 VSS 749 ICV_10 $T=132020 155040 1 0 $X=131830 $Y=152080
X780 VSS VDD 754 ICV_11 $T=145820 13600 0 0 $X=145630 $Y=13360
X781 VSS VDD 754 ICV_11 $T=145820 19040 0 0 $X=145630 $Y=18800
X782 VSS VDD 207 ICV_11 $T=145820 29920 0 0 $X=145630 $Y=29680
X783 VSS VDD 272 ICV_11 $T=145820 46240 0 0 $X=145630 $Y=46000
X784 VSS VDD 754 ICV_11 $T=145820 51680 0 0 $X=145630 $Y=51440
X785 VSS VDD 754 ICV_11 $T=145820 57120 0 0 $X=145630 $Y=56880
X786 VSS VDD 140 ICV_11 $T=145820 84320 0 0 $X=145630 $Y=84080
X787 VSS VDD 140 ICV_11 $T=145820 144160 0 0 $X=145630 $Y=143920
X788 VSS VDD PAR_IN6<13> 59 VDD 78 VSS sky130_fd_sc_hd__and2_4 $T=7820 89760 0 0 $X=7630 $Y=89520
X789 VSS VDD PAR_IN6<29> 59 VDD 79 VSS sky130_fd_sc_hd__and2_4 $T=8280 111520 1 0 $X=8090 $Y=108560
X790 VSS VDD PAR_IN5<12> 67 VDD 87 VSS sky130_fd_sc_hd__and2_4 $T=8280 133280 1 0 $X=8090 $Y=130320
X791 VSS VDD PAR_IN2<25> 66 VDD 106 VSS sky130_fd_sc_hd__and2_4 $T=11500 155040 1 0 $X=11310 $Y=152080
X792 VSS VDD PAR_IN6<25> 103 VDD 111 VSS sky130_fd_sc_hd__and2_4 $T=12420 144160 1 0 $X=12230 $Y=141200
X793 VSS VDD PAR_IN5<4> 67 VDD 112 VSS sky130_fd_sc_hd__and2_4 $T=12880 19040 1 0 $X=12690 $Y=16080
X794 VSS VDD PAR_IN5<29> 89 VDD 114 VSS sky130_fd_sc_hd__and2_4 $T=12880 84320 1 0 $X=12690 $Y=81360
X795 VSS VDD 72 115 VDD 64 VSS sky130_fd_sc_hd__and2_4 $T=16100 46240 0 0 $X=15910 $Y=46000
X796 VSS VDD PAR_IN5<15> 127 VDD 148 VSS sky130_fd_sc_hd__and2_4 $T=20240 122400 0 0 $X=20050 $Y=122160
X797 VSS VDD PAR_IN5<13> 89 VDD 150 VSS sky130_fd_sc_hd__and2_4 $T=22080 29920 0 0 $X=21890 $Y=29680
X798 VSS VDD PAR_IN5<21> 89 VDD 176 VSS sky130_fd_sc_hd__and2_4 $T=23920 13600 0 0 $X=23730 $Y=13360
X799 VSS VDD PAR_IN5<25> 140 VDD 197 VSS sky130_fd_sc_hd__and2_4 $T=28520 155040 1 0 $X=28330 $Y=152080
X800 VSS VDD PAR_IN3<20> 228 VDD 231 VSS sky130_fd_sc_hd__and2_4 $T=40020 13600 0 0 $X=39830 $Y=13360
X801 VSS VDD PAR_IN6<26> 264 VDD 260 VSS sky130_fd_sc_hd__and2_4 $T=48760 19040 0 0 $X=48570 $Y=18800
X802 VSS VDD PAR_IN2<5> 272 VDD 273 VSS sky130_fd_sc_hd__and2_4 $T=49680 68000 1 0 $X=49490 $Y=65040
X803 VSS VDD PAR_IN2<4> 258 VDD 249 VSS sky130_fd_sc_hd__and2_4 $T=49680 138720 1 0 $X=49490 $Y=135760
X804 VSS VDD PAR_IN2<24> 258 VDD 314 VSS sky130_fd_sc_hd__and2_4 $T=54280 149600 1 0 $X=54090 $Y=146640
X805 VSS VDD PAR_IN7<6> 286 VDD 333 VSS sky130_fd_sc_hd__and2_4 $T=57500 78880 1 0 $X=57310 $Y=75920
X806 VSS VDD PAR_IN2<16> 258 VDD 338 VSS sky130_fd_sc_hd__and2_4 $T=58420 106080 1 0 $X=58230 $Y=103120
X807 VSS VDD PAR_IN8<20> 348 VDD 332 VSS sky130_fd_sc_hd__and2_4 $T=63020 35360 0 0 $X=62830 $Y=35120
X808 VSS VDD PAR_IN7<14> 285 VDD 366 VSS sky130_fd_sc_hd__and2_4 $T=63020 106080 0 0 $X=62830 $Y=105840
X809 VSS VDD PAR_IN4<26> 343 VDD 370 VSS sky130_fd_sc_hd__and2_4 $T=63480 116960 0 0 $X=63290 $Y=116720
X810 VSS VDD PAR_IN2<11> 272 VDD 398 VSS sky130_fd_sc_hd__and2_4 $T=66240 19040 1 0 $X=66050 $Y=16080
X811 VSS VDD PAR_IN2<21> 272 VDD 420 VSS sky130_fd_sc_hd__and2_4 $T=78200 19040 0 0 $X=78010 $Y=18800
X812 VSS VDD PAR_IN2<29> 336 VDD 421 VSS sky130_fd_sc_hd__and2_4 $T=93380 46240 1 0 $X=93190 $Y=43280
X813 VSS VDD PAR_IN4<15> 560 VDD 537 VSS sky130_fd_sc_hd__and2_4 $T=97060 95200 0 0 $X=96870 $Y=94960
X814 VSS VDD PAR_IN6<10> 264 VDD 611 VSS sky130_fd_sc_hd__and2_4 $T=105800 29920 1 0 $X=105610 $Y=26960
X815 VSS VDD PAR_IN5<6> 604 VDD 465 VSS sky130_fd_sc_hd__and2_4 $T=105800 68000 1 0 $X=105610 $Y=65040
X816 VSS VDD PAR_IN2<17> 66 VDD 581 VSS sky130_fd_sc_hd__and2_4 $T=107180 51680 0 0 $X=106990 $Y=51440
X817 VSS VDD PAR_IN6<12> 103 VDD 644 VSS sky130_fd_sc_hd__and2_4 $T=109480 144160 0 0 $X=109290 $Y=143920
X818 VSS VDD PAR_IN6<17> 643 VDD 593 VSS sky130_fd_sc_hd__and2_4 $T=110860 13600 0 0 $X=110670 $Y=13360
X819 VSS VDD PAR_IN5<23> 563 VDD 652 VSS sky130_fd_sc_hd__and2_4 $T=112700 149600 1 0 $X=112510 $Y=146640
X820 VSS VDD PAR_IN6<3> 643 VDD 657 VSS sky130_fd_sc_hd__and2_4 $T=113160 19040 1 0 $X=112970 $Y=16080
X821 VSS VDD PAR_IN6<1> 672 VDD 670 VSS sky130_fd_sc_hd__and2_4 $T=119140 127840 0 0 $X=118950 $Y=127600
X822 VSS VDD PAR_IN6<19> 437 VDD 688 VSS sky130_fd_sc_hd__and2_4 $T=119140 155040 1 0 $X=118950 $Y=152080
X823 VSS VDD PAR_IN6<16> 672 VDD 699 VSS sky130_fd_sc_hd__and2_4 $T=120060 116960 1 0 $X=119870 $Y=114000
X824 VSS VDD PAR_IN4<9> 602 VDD 441 VSS sky130_fd_sc_hd__and2_4 $T=120060 149600 1 0 $X=119870 $Y=146640
X825 VSS VDD PAR_IN6<18> 625 VDD 701 VSS sky130_fd_sc_hd__and2_4 $T=120520 144160 1 0 $X=120330 $Y=141200
X826 VSS VDD PAR_IN4<6> 602 VDD 704 VSS sky130_fd_sc_hd__and2_4 $T=120980 116960 0 0 $X=120790 $Y=116720
X827 VSS VDD PAR_IN2<3> 290 VDD 615 VSS sky130_fd_sc_hd__and2_4 $T=122360 57120 1 0 $X=122170 $Y=54160
X828 VSS VDD PAR_IN6<31> 643 VDD 715 VSS sky130_fd_sc_hd__and2_4 $T=123740 19040 1 0 $X=123550 $Y=16080
X829 VSS VDD PAR_IN5<16> 67 VDD 709 VSS sky130_fd_sc_hd__and2_4 $T=128340 13600 0 0 $X=128150 $Y=13360
X830 VSS VDD PAR_IN8<18> 329 VDD 765 VSS sky130_fd_sc_hd__and2_4 $T=133400 57120 1 0 $X=133210 $Y=54160
X831 VSS VDD PAR_IN2<28> 395 VDD 774 VSS sky130_fd_sc_hd__and2_4 $T=134780 116960 0 0 $X=134590 $Y=116720
X832 VSS VDD PAR_IN4<30> 754 VDD 776 VSS sky130_fd_sc_hd__and2_4 $T=137080 46240 0 0 $X=136890 $Y=46000
X833 VSS VDD PAR_IN6<23> 643 VDD 749 VSS sky130_fd_sc_hd__and2_4 $T=138000 155040 1 0 $X=137810 $Y=152080
X834 VSS VDD PAR_IN8<30> 329 VDD 725 VSS sky130_fd_sc_hd__and2_4 $T=138920 84320 0 0 $X=138730 $Y=84080
X835 VSS VDD PAR_IN5<24> 140 VDD 627 VSS sky130_fd_sc_hd__and2_4 $T=143980 149600 1 0 $X=143790 $Y=146640
X836 VSS VDD PAR_IN2<23> 272 VDD 792 VSS sky130_fd_sc_hd__and2_4 $T=144900 78880 1 0 $X=144710 $Y=75920
X837 VSS VDD ICV_12 $T=17940 13600 1 0 $X=17750 $Y=10640
X838 VSS VDD ICV_12 $T=17940 116960 1 0 $X=17750 $Y=114000
X839 VSS VDD ICV_12 $T=17940 155040 0 0 $X=17750 $Y=154800
X840 VSS VDD ICV_12 $T=46000 62560 1 0 $X=45810 $Y=59600
X841 VSS VDD ICV_12 $T=46000 84320 1 0 $X=45810 $Y=81360
X842 VSS VDD ICV_12 $T=74060 149600 1 0 $X=73870 $Y=146640
X843 VSS VDD ICV_12 $T=102120 51680 1 0 $X=101930 $Y=48720
X844 VSS VDD ICV_12 $T=130180 138720 1 0 $X=129990 $Y=135760
X845 VSS VDD ICV_12 $T=143980 62560 0 0 $X=143790 $Y=62320
X846 VSS VDD ICV_12 $T=143980 78880 0 0 $X=143790 $Y=78640
X847 VSS VDD 49 ICV_13 $T=7820 24480 0 0 $X=7630 $Y=24240
X848 VSS VDD 58 ICV_13 $T=7820 78880 1 0 $X=7630 $Y=75920
X849 VSS VDD 60 ICV_13 $T=7820 106080 1 0 $X=7630 $Y=103120
X850 VSS VDD 91 ICV_13 $T=11500 116960 1 0 $X=11310 $Y=114000
X851 VSS VDD 102 ICV_13 $T=12420 133280 1 0 $X=12230 $Y=130320
X852 VSS VDD 105 ICV_13 $T=13340 24480 1 0 $X=13150 $Y=21520
X853 VSS VDD 203 ICV_13 $T=35880 116960 1 0 $X=35690 $Y=114000
X854 VSS VDD 204 ICV_13 $T=37260 35360 1 0 $X=37070 $Y=32400
X855 VSS VDD 165 ICV_13 $T=38180 29920 1 0 $X=37990 $Y=26960
X856 VSS VDD 232 ICV_13 $T=40480 68000 1 0 $X=40290 $Y=65040
X857 VSS VDD 143 ICV_13 $T=40940 57120 1 0 $X=40750 $Y=54160
X858 VSS VDD 229 ICV_13 $T=43700 84320 0 0 $X=43510 $Y=84080
X859 VSS VDD PAR_IN3<20> ICV_13 $T=44160 13600 0 0 $X=43970 $Y=13360
X860 VSS VDD 264 ICV_13 $T=49220 19040 1 0 $X=49030 $Y=16080
X861 VSS VDD SAMPLE_COUNT<1> ICV_13 $T=51520 29920 1 0 $X=51330 $Y=26960
X862 VSS VDD 203 ICV_13 $T=53360 144160 1 0 $X=53170 $Y=141200
X863 VSS VDD 228 ICV_13 $T=53820 95200 0 0 $X=53630 $Y=94960
X864 VSS VDD 283 ICV_13 $T=53820 138720 1 0 $X=53630 $Y=135760
X865 VSS VDD 102 ICV_13 $T=66700 155040 1 0 $X=66510 $Y=152080
X866 VSS VDD 389 ICV_13 $T=67620 149600 1 0 $X=67430 $Y=146640
X867 VSS VDD 394 ICV_13 $T=68080 73440 1 0 $X=67890 $Y=70480
X868 VSS VDD 314 ICV_13 $T=69460 133280 1 0 $X=69270 $Y=130320
X869 VSS VDD 391 ICV_13 $T=72680 46240 0 0 $X=72490 $Y=46000
X870 VSS VDD 436 ICV_13 $T=77280 84320 1 0 $X=77090 $Y=81360
X871 VSS VDD 401 ICV_13 $T=78200 13600 1 0 $X=78010 $Y=10640
X872 VSS VDD 348 ICV_13 $T=78200 62560 0 0 $X=78010 $Y=62320
X873 VSS VDD 386 ICV_13 $T=80040 46240 0 0 $X=79850 $Y=46000
X874 VSS VDD 453 ICV_13 $T=81420 138720 0 0 $X=81230 $Y=138480
X875 VSS VDD 456 ICV_13 $T=88320 89760 1 0 $X=88130 $Y=86800
X876 VSS VDD 513 ICV_13 $T=90160 155040 1 0 $X=89970 $Y=152080
X877 VSS VDD 303 ICV_13 $T=91080 51680 0 0 $X=90890 $Y=51440
X878 VSS VDD 304 ICV_13 $T=91080 144160 1 0 $X=90890 $Y=141200
X879 VSS VDD 546 ICV_13 $T=95680 51680 1 0 $X=95490 $Y=48720
X880 VSS VDD 549 ICV_13 $T=96140 35360 1 0 $X=95950 $Y=32400
X881 VSS VDD 559 ICV_13 $T=97520 46240 1 0 $X=97330 $Y=43280
X882 VSS VDD 517 ICV_13 $T=97980 73440 0 0 $X=97790 $Y=73200
X883 VSS VDD 556 ICV_13 $T=98440 89760 0 0 $X=98250 $Y=89520
X884 VSS VDD 66 ICV_13 $T=105340 149600 1 0 $X=105150 $Y=146640
X885 VSS VDD 602 ICV_13 $T=105800 138720 0 0 $X=105610 $Y=138480
X886 VSS VDD 468 ICV_13 $T=109020 78880 1 0 $X=108830 $Y=75920
X887 VSS VDD 637 ICV_13 $T=109940 111520 1 0 $X=109750 $Y=108560
X888 VSS VDD 66 ICV_13 $T=110400 57120 1 0 $X=110210 $Y=54160
X889 VSS VDD 672 ICV_13 $T=118220 127840 1 0 $X=118030 $Y=124880
X890 VSS VDD 677 ICV_13 $T=118680 138720 1 0 $X=118490 $Y=135760
X891 VSS VDD 620 ICV_13 $T=120060 24480 1 0 $X=119870 $Y=21520
X892 VSS VDD 127 ICV_13 $T=120980 13600 1 0 $X=120790 $Y=10640
X893 VSS VDD 374 ICV_13 $T=122820 100640 1 0 $X=122630 $Y=97680
X894 VSS VDD PAR_IN8<0> ICV_13 $T=123280 155040 1 0 $X=123090 $Y=152080
X895 VSS VDD PAR_IN2<3> ICV_13 $T=125580 51680 0 0 $X=125390 $Y=51440
X896 VSS VDD 688 ICV_13 $T=125580 73440 1 0 $X=125390 $Y=70480
X897 VSS VDD 374 ICV_13 $T=125580 73440 0 0 $X=125390 $Y=73200
X898 VSS VDD 643 ICV_13 $T=136160 13600 0 0 $X=135970 $Y=13360
X899 VSS VDD 765 ICV_13 $T=137540 62560 0 0 $X=137350 $Y=62320
X900 VSS VDD PAR_IN2<28> ICV_13 $T=138920 116960 0 0 $X=138730 $Y=116720
X901 VSS VDD 653 ICV_13 $T=139380 40800 1 0 $X=139190 $Y=37840
X902 VSS VDD 792 ICV_13 $T=141220 68000 1 0 $X=141030 $Y=65040
X903 VSS VDD 329 ICV_13 $T=142600 111520 1 0 $X=142410 $Y=108560
X904 VSS VDD 285 ICV_13 $T=143520 100640 1 0 $X=143330 $Y=97680
X905 VSS VDD PAR_IN5<2> 271 391 ICV_14 $T=66700 46240 1 0 $X=66510 $Y=43280
X906 VSS VDD PAR_IN6<7> 437 486 ICV_14 $T=81420 155040 1 0 $X=81230 $Y=152080
X907 VSS VDD PAR_IN6<27> 643 767 ICV_14 $T=133400 19040 1 0 $X=133210 $Y=16080
X908 VSS VDD PAR_IN7<20> 617 371 ICV_14 $T=141680 29920 1 0 $X=141490 $Y=26960
X909 VSS VDD PAR_IN7<2> 285 738 ICV_14 $T=142600 106080 1 0 $X=142410 $Y=103120
X910 VSS VDD PAR_IN8<26> 329 668 ICV_14 $T=142600 116960 1 0 $X=142410 $Y=114000
X911 VSS VDD PAR_IN4<22> 754 621 ICV_14 $T=143060 24480 1 0 $X=142870 $Y=21520
X912 VSS VDD PAR_IN2<27> 272 740 ICV_14 $T=143060 51680 1 0 $X=142870 $Y=48720
X913 VSS VDD PAR_IN4<18> 754 762 ICV_14 $T=143520 19040 1 0 $X=143330 $Y=16080
X914 VSS VDD PAR_IN4<2> 754 781 ICV_14 $T=143520 62560 1 0 $X=143330 $Y=59600
X915 VSS VDD PAR_IN5<28> 140 796 ICV_14 $T=143520 89760 1 0 $X=143330 $Y=86800
X916 VSS VDD SAMPLE_COUNT<2> ICV_15 $T=7820 40800 1 0 $X=7630 $Y=37840
X917 VSS VDD 81 ICV_15 $T=14260 133280 0 0 $X=14070 $Y=133040
X918 VSS VDD 4 ICV_15 $T=22080 24480 0 0 $X=21890 $Y=24240
X919 VSS VDD 97 ICV_15 $T=26220 95200 1 0 $X=26030 $Y=92240
X920 VSS VDD 69 ICV_15 $T=31280 57120 0 0 $X=31090 $Y=56880
X921 VSS VDD 165 ICV_15 $T=31280 106080 0 0 $X=31090 $Y=105840
X922 VSS VDD 286 ICV_15 $T=52440 73440 1 0 $X=52250 $Y=70480
X923 VSS VDD 248 ICV_15 $T=52440 111520 0 0 $X=52250 $Y=111280
X924 VSS VDD 290 ICV_15 $T=54740 13600 1 0 $X=54550 $Y=10640
X925 VSS VDD 348 ICV_15 $T=62560 40800 1 0 $X=62370 $Y=37840
X926 VSS VDD 285 ICV_15 $T=62560 106080 1 0 $X=62370 $Y=103120
X927 VSS VDD 271 ICV_15 $T=68540 40800 1 0 $X=68350 $Y=37840
X928 VSS VDD 434 ICV_15 $T=77280 73440 1 0 $X=77090 $Y=70480
X929 VSS VDD 459 ICV_15 $T=83720 100640 0 0 $X=83530 $Y=100400
X930 VSS VDD 621 ICV_15 $T=107640 106080 1 0 $X=107450 $Y=103120
X931 VSS VDD 643 ICV_15 $T=110860 13600 1 0 $X=110670 $Y=10640
X932 VSS VDD 563 ICV_15 $T=112700 144160 1 0 $X=112510 $Y=141200
X933 VSS VDD 137 ICV_15 $T=115460 62560 0 0 $X=115270 $Y=62320
X934 VSS VDD 655 ICV_15 $T=115460 73440 0 0 $X=115270 $Y=73200
X935 VSS VDD 620 ICV_15 $T=115460 89760 0 0 $X=115270 $Y=89520
X936 VSS VDD PAR_IN6<16> ICV_15 $T=125580 111520 0 0 $X=125390 $Y=111280
X937 VSS VDD PAR_IN4<28> ICV_15 $T=132480 116960 0 0 $X=132290 $Y=116720
X938 VSS VDD 329 ICV_15 $T=138920 84320 1 0 $X=138730 $Y=81360
X939 VSS VDD PAR_IN4<18> ICV_15 $T=143520 13600 0 0 $X=143330 $Y=13360
X940 VSS VDD PAR_IN4<2> ICV_15 $T=143520 57120 0 0 $X=143330 $Y=56880
X941 VSS VDD RESET ICV_16 $T=7820 29920 1 0 $X=7630 $Y=26960
X942 VSS VDD 55 ICV_16 $T=7820 35360 1 0 $X=7630 $Y=32400
X943 VSS VDD 66 ICV_16 $T=8280 122400 1 0 $X=8090 $Y=119440
X944 VSS VDD 67 ICV_16 $T=8280 127840 1 0 $X=8090 $Y=124880
X945 VSS VDD PAR_IN5<12> ICV_16 $T=8280 127840 0 0 $X=8090 $Y=127600
X946 VSS VDD 80 ICV_16 $T=9660 144160 1 0 $X=9470 $Y=141200
X947 VSS VDD 5 ICV_16 $T=16560 51680 1 0 $X=16370 $Y=48720
X948 VSS VDD 64 ICV_16 $T=17020 35360 1 0 $X=16830 $Y=32400
X949 VSS VDD CLK ICV_16 $T=20700 68000 0 0 $X=20510 $Y=67760
X950 VSS VDD 56 ICV_16 $T=21160 57120 1 0 $X=20970 $Y=54160
X951 VSS VDD 133 ICV_16 $T=21160 89760 0 0 $X=20970 $Y=89520
X952 VSS VDD 69 ICV_16 $T=24840 46240 1 0 $X=24650 $Y=43280
X953 VSS VDD 116 ICV_16 $T=27600 84320 1 0 $X=27410 $Y=81360
X954 VSS VDD 81 ICV_16 $T=28520 122400 0 0 $X=28330 $Y=122160
X955 VSS VDD 165 ICV_16 $T=28980 19040 0 0 $X=28790 $Y=18800
X956 VSS VDD 193 ICV_16 $T=30360 78880 0 0 $X=30170 $Y=78640
X957 VSS VDD 191 ICV_16 $T=30820 40800 0 0 $X=30630 $Y=40560
X958 VSS VDD COUNT<5> ICV_16 $T=30820 68000 0 0 $X=30630 $Y=67760
X959 VSS VDD 30 ICV_16 $T=30820 95200 0 0 $X=30630 $Y=94960
X960 VSS VDD 183 ICV_16 $T=30820 100640 0 0 $X=30630 $Y=100400
X961 VSS VDD PAR_IN5<25> ICV_16 $T=30820 149600 0 0 $X=30630 $Y=149360
X962 VSS VDD 11 ICV_16 $T=34500 84320 1 0 $X=34310 $Y=81360
X963 VSS VDD 193 ICV_16 $T=34960 84320 0 0 $X=34770 $Y=84080
X964 VSS VDD 13 ICV_16 $T=34960 95200 1 0 $X=34770 $Y=92240
X965 VSS VDD COUNT<0> ICV_16 $T=37260 68000 0 0 $X=37070 $Y=67760
X966 VSS VDD PAR_IN8<8> ICV_16 $T=37260 138720 0 0 $X=37070 $Y=138480
X967 VSS VDD SAMPLE_COUNT<3> ICV_16 $T=37720 68000 1 0 $X=37530 $Y=65040
X968 VSS VDD SAMPLE_COUNT<3> ICV_16 $T=40020 40800 0 0 $X=39830 $Y=40560
X969 VSS VDD 222 ICV_16 $T=40940 89760 1 0 $X=40750 $Y=86800
X970 VSS VDD 4 ICV_16 $T=41400 51680 0 0 $X=41210 $Y=51440
X971 VSS VDD 229 ICV_16 $T=42320 111520 0 0 $X=42130 $Y=111280
X972 VSS VDD 193 ICV_16 $T=43700 73440 0 0 $X=43510 $Y=73200
X973 VSS VDD 237 ICV_16 $T=45080 122400 1 0 $X=44890 $Y=119440
X974 VSS VDD 218 ICV_16 $T=48300 127840 0 0 $X=48110 $Y=127600
X975 VSS VDD 70 ICV_16 $T=49680 73440 1 0 $X=49490 $Y=70480
X976 VSS VDD COUNT<1> ICV_16 $T=51060 89760 0 0 $X=50870 $Y=89520
X977 VSS VDD 265 ICV_16 $T=51980 40800 0 0 $X=51790 $Y=40560
X978 VSS VDD 211 ICV_16 $T=56120 51680 1 0 $X=55930 $Y=48720
X979 VSS VDD 319 ICV_16 $T=57040 106080 0 0 $X=56850 $Y=105840
X980 VSS VDD PAR_IN2<7> ICV_16 $T=58880 24480 0 0 $X=58690 $Y=24240
X981 VSS VDD SAMPLE_COUNT<3> ICV_16 $T=58880 46240 0 0 $X=58690 $Y=46000
X982 VSS VDD 239 ICV_16 $T=63020 40800 0 0 $X=62830 $Y=40560
X983 VSS VDD 300 ICV_16 $T=63020 51680 1 0 $X=62830 $Y=48720
X984 VSS VDD COUNT<1> ICV_16 $T=73600 95200 0 0 $X=73410 $Y=94960
X985 VSS VDD 433 ICV_16 $T=77280 57120 1 0 $X=77090 $Y=54160
X986 VSS VDD PAR_IN1<20> ICV_16 $T=80040 13600 0 0 $X=79850 $Y=13360
X987 VSS VDD 426 ICV_16 $T=82340 40800 1 0 $X=82150 $Y=37840
X988 VSS VDD 271 ICV_16 $T=85100 57120 1 0 $X=84910 $Y=54160
X989 VSS VDD 202 ICV_16 $T=85100 95200 0 0 $X=84910 $Y=94960
X990 VSS VDD PAR_IN1<11> ICV_16 $T=86480 78880 0 0 $X=86290 $Y=78640
X991 VSS VDD PAR_IN7<21> ICV_16 $T=86940 24480 0 0 $X=86750 $Y=24240
X992 VSS VDD 511 ICV_16 $T=89240 62560 1 0 $X=89050 $Y=59600
X993 VSS VDD PAR_IN3<22> ICV_16 $T=91540 100640 1 0 $X=91350 $Y=97680
X994 VSS VDD 388 ICV_16 $T=92000 133280 0 0 $X=91810 $Y=133040
X995 VSS VDD 181 ICV_16 $T=94760 122400 0 0 $X=94570 $Y=122160
X996 VSS VDD PAR_IN5<3> ICV_16 $T=97520 149600 0 0 $X=97330 $Y=149360
X997 VSS VDD 228 ICV_16 $T=97980 68000 0 0 $X=97790 $Y=67760
X998 VSS VDD PAR_IN1<29> ICV_16 $T=103500 29920 0 0 $X=103310 $Y=29680
X999 VSS VDD PAR_IN1<5> ICV_16 $T=104880 78880 0 0 $X=104690 $Y=78640
X1000 VSS VDD 595 ICV_16 $T=105340 51680 1 0 $X=105150 $Y=48720
X1001 VSS VDD 392 ICV_16 $T=106260 35360 1 0 $X=106070 $Y=32400
X1002 VSS VDD 103 ICV_16 $T=109480 144160 1 0 $X=109290 $Y=141200
X1003 VSS VDD PAR_IN4<10> ICV_16 $T=114540 116960 0 0 $X=114350 $Y=116720
X1004 VSS VDD 631 ICV_16 $T=115000 24480 0 0 $X=114810 $Y=24240
X1005 VSS VDD PAR_IN7<10> ICV_16 $T=115000 95200 0 0 $X=114810 $Y=94960
X1006 VSS VDD 271 ICV_16 $T=119140 46240 0 0 $X=118950 $Y=46000
X1007 VSS VDD 652 ICV_16 $T=122820 84320 0 0 $X=122630 $Y=84080
X1008 VSS VDD PAR_IN5<9> ICV_16 $T=123280 24480 0 0 $X=123090 $Y=24240
X1009 VSS VDD 699 ICV_16 $T=125120 111520 1 0 $X=124930 $Y=108560
X1010 VSS VDD 672 ICV_16 $T=126960 122400 1 0 $X=126770 $Y=119440
X1011 VSS VDD 730 ICV_16 $T=128800 62560 1 0 $X=128610 $Y=59600
X1012 VSS VDD 752 ICV_16 $T=133400 122400 0 0 $X=133210 $Y=122160
X1013 VSS VDD 343 ICV_16 $T=133860 46240 0 0 $X=133670 $Y=46000
X1014 VSS VDD 754 ICV_16 $T=137080 51680 1 0 $X=136890 $Y=48720
X1015 VSS VDD 617 ICV_16 $T=138460 138720 1 0 $X=138270 $Y=135760
X1016 VSS VDD PAR_IN6<2> ICV_16 $T=139840 51680 1 0 $X=139650 $Y=48720
X1017 VSS VDD PAR_IN8<5> ICV_16 $T=140300 89760 1 0 $X=140110 $Y=86800
X1018 VSS VDD PAR_IN4<22> ICV_16 $T=143060 19040 0 0 $X=142870 $Y=18800
X1019 VSS VDD 653 ICV_16 $T=143060 95200 0 0 $X=142870 $Y=94960
X1020 VSS VDD PAR_IN7<2> ICV_16 $T=143060 100640 0 0 $X=142870 $Y=100400
X1021 VSS VDD PAR_IN2<0> ICV_16 $T=143060 133280 0 0 $X=142870 $Y=133040
X1022 VSS VDD 85 ICV_17 $T=11500 122400 1 0 $X=11310 $Y=119440
X1023 VSS VDD 81 ICV_17 $T=17020 149600 0 0 $X=16830 $Y=149360
X1024 VSS VDD 113 ICV_17 $T=24380 62560 0 0 $X=24190 $Y=62320
X1025 VSS VDD 164 ICV_17 $T=24380 155040 1 0 $X=24190 $Y=152080
X1026 VSS VDD 235 ICV_17 $T=43700 138720 1 0 $X=43510 $Y=135760
X1027 VSS VDD 246 ICV_17 $T=44160 89760 1 0 $X=43970 $Y=86800
X1028 VSS VDD SAMPLE_COUNT<1> ICV_17 $T=49220 24480 0 0 $X=49030 $Y=24240
X1029 VSS VDD 268 ICV_17 $T=55200 40800 1 0 $X=55010 $Y=37840
X1030 VSS VDD 178 ICV_17 $T=55660 84320 0 0 $X=55470 $Y=84080
X1031 VSS VDD 262 ICV_17 $T=56120 133280 0 0 $X=55930 $Y=133040
X1032 VSS VDD 274 ICV_17 $T=57500 116960 0 0 $X=57310 $Y=116720
X1033 VSS VDD PAR_IN4<26> ICV_17 $T=67620 116960 0 0 $X=67430 $Y=116720
X1034 VSS VDD PAR_IN5<20> ICV_17 $T=68080 35360 1 0 $X=67890 $Y=32400
X1035 VSS VDD 398 ICV_17 $T=70380 19040 1 0 $X=70190 $Y=16080
X1036 VSS VDD 412 ICV_17 $T=71760 127840 1 0 $X=71570 $Y=124880
X1037 VSS VDD PAR_IN1<13> ICV_17 $T=72680 51680 0 0 $X=72490 $Y=51440
X1038 VSS VDD 482 ICV_17 $T=85560 84320 0 0 $X=85370 $Y=84080
X1039 VSS VDD 91 ICV_17 $T=99820 57120 1 0 $X=99630 $Y=54160
X1040 VSS VDD 148 ICV_17 $T=100280 122400 1 0 $X=100090 $Y=119440
X1041 VSS VDD PAR_IN6<5> ICV_17 $T=101660 155040 0 0 $X=101470 $Y=154800
X1042 VSS VDD 615 ICV_17 $T=109940 57120 0 0 $X=109750 $Y=56880
X1043 VSS VDD 619 ICV_17 $T=109940 68000 1 0 $X=109750 $Y=65040
X1044 VSS VDD 282 ICV_17 $T=109940 78880 0 0 $X=109750 $Y=78640
X1045 VSS VDD 271 ICV_17 $T=113620 57120 0 0 $X=113430 $Y=56880
X1046 VSS VDD 604 ICV_17 $T=121440 89760 0 0 $X=121250 $Y=89520
X1047 VSS VDD 602 ICV_17 $T=124200 116960 1 0 $X=124010 $Y=114000
X1048 VSS VDD 395 ICV_17 $T=127880 84320 1 0 $X=127690 $Y=81360
X1049 VSS VDD 725 ICV_17 $T=127880 89760 1 0 $X=127690 $Y=86800
X1050 VSS VDD 285 ICV_17 $T=132480 73440 0 0 $X=132290 $Y=73200
X1051 VSS VDD 546 ICV_17 $T=138000 24480 0 0 $X=137810 $Y=24240
X1052 VSS VDD 338 ICV_17 $T=138460 116960 1 0 $X=138270 $Y=114000
X1053 VSS VDD PAR_IN6<24> ICV_17 $T=142140 122400 0 0 $X=141950 $Y=122160
X1054 VSS VDD 64 ICV_18 $T=6900 51680 1 0 $X=6710 $Y=48720
X1055 VSS VDD 5 ICV_18 $T=6900 57120 1 0 $X=6710 $Y=54160
X1056 VSS VDD INTERNAL_FINISH ICV_18 $T=6900 68000 0 0 $X=6710 $Y=67760
X1057 VSS VDD 12 ICV_18 $T=11040 89760 0 0 $X=10850 $Y=89520
X1058 VSS VDD 113 ICV_18 $T=14260 78880 1 0 $X=14070 $Y=75920
X1059 VSS VDD 137 ICV_18 $T=20240 111520 1 0 $X=20050 $Y=108560
X1060 VSS VDD 138 ICV_18 $T=20240 116960 1 0 $X=20050 $Y=114000
X1061 VSS VDD 150 ICV_18 $T=23920 73440 1 0 $X=23730 $Y=70480
X1062 VSS VDD 164 ICV_18 $T=24380 138720 1 0 $X=24190 $Y=135760
X1063 VSS VDD PAR_IN1<26> ICV_18 $T=30360 127840 0 0 $X=30170 $Y=127600
X1064 VSS VDD 12 ICV_18 $T=31280 89760 1 0 $X=31090 $Y=86800
X1065 VSS VDD 206 ICV_18 $T=32660 133280 1 0 $X=32470 $Y=130320
X1066 VSS VDD 13 ICV_18 $T=37720 95200 0 0 $X=37530 $Y=94960
X1067 VSS VDD 143 ICV_18 $T=44620 40800 1 0 $X=44430 $Y=37840
X1068 VSS VDD PAR_IN6<26> ICV_18 $T=45540 19040 0 0 $X=45350 $Y=18800
X1069 VSS VDD 343 ICV_18 $T=62100 122400 1 0 $X=61910 $Y=119440
X1070 VSS VDD PAR_IN3<11> ICV_18 $T=65780 19040 0 0 $X=65590 $Y=18800
X1071 VSS VDD 374 ICV_18 $T=67620 89760 1 0 $X=67430 $Y=86800
X1072 VSS VDD 406 ICV_18 $T=68540 138720 1 0 $X=68350 $Y=135760
X1073 VSS VDD 373 ICV_18 $T=77740 106080 0 0 $X=77550 $Y=105840
X1074 VSS VDD 341 ICV_18 $T=80040 122400 1 0 $X=79850 $Y=119440
X1075 VSS VDD 476 ICV_18 $T=81420 100640 1 0 $X=81230 $Y=97680
X1076 VSS VDD 479 ICV_18 $T=81880 68000 1 0 $X=81690 $Y=65040
X1077 VSS VDD 413 ICV_18 $T=86480 40800 0 0 $X=86290 $Y=40560
X1078 VSS VDD 457 ICV_18 $T=86480 46240 0 0 $X=86290 $Y=46000
X1079 VSS VDD 502 ICV_18 $T=86480 116960 0 0 $X=86290 $Y=116720
X1080 VSS VDD 529 ICV_18 $T=90620 122400 1 0 $X=90430 $Y=119440
X1081 VSS VDD PAR_IN6<14> ICV_18 $T=92000 46240 0 0 $X=91810 $Y=46000
X1082 VSS VDD 550 ICV_18 $T=94760 57120 1 0 $X=94570 $Y=54160
X1083 VSS VDD PAR_IN7<15> ICV_18 $T=95220 127840 0 0 $X=95030 $Y=127600
X1084 VSS VDD 480 ICV_18 $T=96600 116960 1 0 $X=96410 $Y=114000
X1085 VSS VDD 585 ICV_18 $T=100740 68000 1 0 $X=100550 $Y=65040
X1086 VSS VDD 620 ICV_18 $T=106260 100640 1 0 $X=106070 $Y=97680
X1087 VSS VDD 264 ICV_18 $T=110860 35360 1 0 $X=110670 $Y=32400
X1088 VSS VDD 659 ICV_18 $T=114080 68000 0 0 $X=113890 $Y=67760
X1089 VSS VDD 164 ICV_18 $T=116840 57120 1 0 $X=116650 $Y=54160
X1090 VSS VDD 654 ICV_18 $T=124660 78880 0 0 $X=124470 $Y=78640
X1091 VSS VDD PAR_IN7<24> ICV_18 $T=124660 133280 0 0 $X=124470 $Y=133040
X1092 VSS VDD 546 ICV_18 $T=135700 51680 0 0 $X=135510 $Y=51440
X1093 VSS VDD 781 ICV_18 $T=136620 57120 1 0 $X=136430 $Y=54160
X1094 VSS VDD PAR_IN5<28> ICV_18 $T=142140 84320 0 0 $X=141950 $Y=84080
X1095 VSS VDD 78 77 PAR_IN7<13> VDD 70 VSS sky130_fd_sc_hd__a21o_4 $T=7820 89760 1 0 $X=7630 $Y=86800
X1096 VSS VDD 79 77 PAR_IN7<29> VDD 71 VSS sky130_fd_sc_hd__a21o_4 $T=7820 111520 0 0 $X=7630 $Y=111280
X1097 VSS VDD 81 80 PAR_IN4<25> VDD 93 VSS sky130_fd_sc_hd__a21o_4 $T=10580 149600 0 0 $X=10390 $Y=149360
X1098 VSS VDD 87 102 PAR_IN8<12> VDD 94 VSS sky130_fd_sc_hd__a21o_4 $T=11040 127840 0 0 $X=10850 $Y=127600
X1099 VSS VDD 116 25 97 VDD 108 VSS sky130_fd_sc_hd__a21o_4 $T=21160 89760 1 0 $X=20970 $Y=86800
X1100 VSS VDD 205 SERIAL_OUT 6 VDD 161 VSS sky130_fd_sc_hd__a21o_4 $T=31740 29920 1 0 $X=31550 $Y=26960
X1101 VSS VDD 188 207 PAR_IN8<8> VDD 187 VSS sky130_fd_sc_hd__a21o_4 $T=34960 144160 1 0 $X=34770 $Y=141200
X1102 VSS VDD 249 178 PAR_IN3<4> VDD 238 VSS sky130_fd_sc_hd__a21o_4 $T=42320 144160 0 0 $X=42130 $Y=143920
X1103 VSS VDD 332 336 PAR_IN2<20> VDD 347 VSS sky130_fd_sc_hd__a21o_4 $T=61640 35360 1 0 $X=61450 $Y=32400
X1104 VSS VDD 333 290 PAR_IN2<6> VDD 352 VSS sky130_fd_sc_hd__a21o_4 $T=62100 89760 1 0 $X=61910 $Y=86800
X1105 VSS VDD 391 373 PAR_IN8<2> VDD 381 VSS sky130_fd_sc_hd__a21o_4 $T=66240 46240 0 0 $X=66050 $Y=46000
X1106 VSS VDD 441 437 PAR_IN6<9> VDD 324 VSS sky130_fd_sc_hd__a21o_4 $T=75900 149600 0 0 $X=75710 $Y=149360
X1107 VSS VDD 457 510 PAR_IN3<14> VDD 446 VSS sky130_fd_sc_hd__a21o_4 $T=89240 51680 1 0 $X=89050 $Y=48720
X1108 VSS VDD 468 431 PAR_IN4<5> VDD 516 VSS sky130_fd_sc_hd__a21o_4 $T=91540 24480 1 0 $X=91350 $Y=21520
X1109 VSS VDD 548 432 PAR_IN8<1> VDD 524 VSS sky130_fd_sc_hd__a21o_4 $T=93840 122400 1 0 $X=93650 $Y=119440
X1110 VSS VDD 559 546 PAR_IN6<14> VDD 429 VSS sky130_fd_sc_hd__a21o_4 $T=95220 46240 0 0 $X=95030 $Y=46000
X1111 VSS VDD 468 431 PAR_IN4<21> VDD 522 VSS sky130_fd_sc_hd__a21o_4 $T=97980 19040 0 0 $X=97790 $Y=18800
X1112 VSS VDD 575 513 PAR_IN7<5> VDD 547 VSS sky130_fd_sc_hd__a21o_4 $T=100280 149600 0 0 $X=100090 $Y=149360
X1113 VSS VDD 493 91 PAR_IN3<15> VDD 591 VSS sky130_fd_sc_hd__a21o_4 $T=103500 127840 0 0 $X=103310 $Y=127600
X1114 VSS VDD 468 431 PAR_IN4<11> VDD 585 VSS sky130_fd_sc_hd__a21o_4 $T=105340 84320 1 0 $X=105150 $Y=81360
X1115 VSS VDD 493 181 PAR_IN4<17> VDD 587 VSS sky130_fd_sc_hd__a21o_4 $T=106720 46240 0 0 $X=106530 $Y=46000
X1116 VSS VDD 624 617 PAR_IN7<22> VDD 571 VSS sky130_fd_sc_hd__a21o_4 $T=107180 111520 0 0 $X=106990 $Y=111280
X1117 VSS VDD 619 137 PAR_IN8<19> VDD 633 VSS sky130_fd_sc_hd__a21o_4 $T=108560 68000 0 0 $X=108370 $Y=67760
X1118 VSS VDD 635 620 PAR_IN5<10> VDD 609 VSS sky130_fd_sc_hd__a21o_4 $T=113160 95200 1 0 $X=112970 $Y=92240
X1119 VSS VDD 593 164 PAR_IN7<17> VDD 578 VSS sky130_fd_sc_hd__a21o_4 $T=113620 24480 1 0 $X=113430 $Y=21520
X1120 VSS VDD 611 286 PAR_IN7<10> VDD 610 VSS sky130_fd_sc_hd__a21o_4 $T=114540 100640 1 0 $X=114350 $Y=97680
X1121 VSS VDD 667 653 PAR_IN4<31> VDD 640 VSS sky130_fd_sc_hd__a21o_4 $T=117300 40800 1 0 $X=117110 $Y=37840
X1122 VSS VDD 657 164 PAR_IN7<3> VDD 588 VSS sky130_fd_sc_hd__a21o_4 $T=119140 51680 0 0 $X=118950 $Y=51440
X1123 VSS VDD 766 77 PAR_IN7<11> VDD 586 VSS sky130_fd_sc_hd__a21o_4 $T=133400 78880 0 0 $X=133210 $Y=78640
X1124 VSS VDD 304 560 PAR_IN4<28> VDD 736 VSS sky130_fd_sc_hd__a21o_4 $T=133400 122400 1 0 $X=133210 $Y=119440
X1125 VSS VDD 740 289 PAR_IN3<27> VDD 772 VSS sky130_fd_sc_hd__a21o_4 $T=136160 46240 1 0 $X=135970 $Y=43280
X1126 VSS VDD 304 560 PAR_IN4<16> VDD 727 VSS sky130_fd_sc_hd__a21o_4 $T=136160 111520 1 0 $X=135970 $Y=108560
X1127 VSS VDD 781 546 PAR_IN6<2> VDD 745 VSS sky130_fd_sc_hd__a21o_4 $T=139840 57120 1 0 $X=139650 $Y=54160
X1128 VSS VDD 792 289 PAR_IN3<23> VDD 746 VSS sky130_fd_sc_hd__a21o_4 $T=141220 73440 1 0 $X=141030 $Y=70480
X1129 VSS VDD 796 207 PAR_IN8<28> VDD 747 VSS sky130_fd_sc_hd__a21o_4 $T=141220 84320 1 0 $X=141030 $Y=81360
X1130 VSS VDD 788 387 PAR_IN3<0> VDD 760 VSS sky130_fd_sc_hd__a21o_4 $T=141680 138720 1 0 $X=141490 $Y=135760
X1131 VSS VDD PAR_IN2<4> 258 ICV_19 $T=49680 133280 0 0 $X=49490 $Y=133040
X1132 VSS VDD 178 304 ICV_19 $T=53360 155040 1 0 $X=53170 $Y=152080
X1133 VSS VDD 16 19 ICV_19 $T=57960 89760 1 0 $X=57770 $Y=86800
X1134 VSS VDD 361 379 ICV_19 $T=64860 106080 1 0 $X=64670 $Y=103120
X1135 VSS VDD 340 301 ICV_19 $T=68540 57120 0 0 $X=68350 $Y=56880
X1136 VSS VDD 469 489 ICV_19 $T=92000 62560 1 0 $X=91810 $Y=59600
X1137 VSS VDD 469 543 ICV_19 $T=96600 35360 0 0 $X=96410 $Y=35120
X1138 VSS VDD PAR_IN6<10> 264 ICV_19 $T=105800 24480 0 0 $X=105610 $Y=24240
X1139 VSS VDD PAR_IN6<18> 625 ICV_19 $T=121440 138720 0 0 $X=121250 $Y=138480
X1140 VSS VDD 677 734 ICV_19 $T=127880 133280 1 0 $X=127690 $Y=130320
X1141 VSS VDD 437 PAR_IN6<11> ICV_19 $T=136160 73440 0 0 $X=135970 $Y=73200
X1142 VSS VDD PAR_IN7<20> 617 ICV_19 $T=141680 24480 0 0 $X=141490 $Y=24240
X1143 VSS VDD ICV_20 $T=6900 13600 1 0 $X=6710 $Y=10640
X1144 VSS VDD ICV_20 $T=6900 155040 0 0 $X=6710 $Y=154800
X1145 VSS VDD ICV_20 $T=20240 155040 0 0 $X=20050 $Y=154800
X1146 VSS VDD ICV_20 $T=22540 116960 1 0 $X=22350 $Y=114000
X1147 VSS VDD ICV_20 $T=29440 62560 1 0 $X=29250 $Y=59600
X1148 VSS VDD ICV_20 $T=33580 40800 1 0 $X=33390 $Y=37840
X1149 VSS VDD ICV_20 $T=34040 62560 0 0 $X=33850 $Y=62320
X1150 VSS VDD ICV_20 $T=34040 100640 1 0 $X=33850 $Y=97680
X1151 VSS VDD ICV_20 $T=35880 24480 1 0 $X=35690 $Y=21520
X1152 VSS VDD ICV_20 $T=37720 24480 0 0 $X=37530 $Y=24240
X1153 VSS VDD ICV_20 $T=54280 100640 1 0 $X=54090 $Y=97680
X1154 VSS VDD ICV_20 $T=94300 138720 0 0 $X=94110 $Y=138480
X1155 VSS VDD ICV_20 $T=118680 95200 1 0 $X=118490 $Y=92240
X1156 VSS VDD ICV_20 $T=137540 127840 1 0 $X=137350 $Y=124880
X1157 VSS VDD ICV_20 $T=138920 122400 1 0 $X=138730 $Y=119440
X1158 VSS VDD ICV_20 $T=141220 155040 1 0 $X=141030 $Y=152080
X1159 VSS VDD 82 97 ICV_21 $T=15180 40800 1 0 $X=14990 $Y=37840
X1160 VSS VDD 98 6 ICV_21 $T=15180 57120 1 0 $X=14990 $Y=54160
X1161 VSS VDD 178 106 ICV_21 $T=28980 144160 0 0 $X=28790 $Y=143920
X1162 VSS VDD SAMPLE_COUNT<0> SAMPLE_COUNT<0> ICV_21 $T=57040 40800 0 0 $X=56850 $Y=40560
X1163 VSS VDD 571 570 ICV_21 $T=99360 106080 1 0 $X=99170 $Y=103120
X1164 VSS VDD 493 181 ICV_21 $T=113160 46240 0 0 $X=112970 $Y=46000
X1165 VSS VDD 687 701 ICV_21 $T=127420 144160 1 0 $X=127230 $Y=141200
X1166 VSS VDD PAR_IN3<23> 289 ICV_21 $T=141220 68000 0 0 $X=141030 $Y=67760
X1167 VSS VDD 72 4 COMPLETE ICV_22 $T=11040 46240 0 0 $X=10850 $Y=46000
X1168 VSS VDD 229 118 219 ICV_22 $T=42320 116960 1 0 $X=42130 $Y=114000
X1169 VSS VDD 351 262 351 ICV_22 $T=63020 138720 0 0 $X=62830 $Y=138480
X1170 VSS VDD 206 303 206 ICV_22 $T=71300 116960 0 0 $X=71110 $Y=116720
X1171 VSS VDD 383 186 186 ICV_22 $T=77740 149600 1 0 $X=77550 $Y=146640
X1172 VSS VDD 348 432 348 ICV_22 $T=84180 35360 0 0 $X=83990 $Y=35120
X1173 VSS VDD 81 468 PAR_IN6<15> ICV_22 $T=92000 95200 0 0 $X=91810 $Y=94960
X1174 VSS VDD 604 127 604 ICV_22 $T=112700 84320 0 0 $X=112510 $Y=84080
X1175 VSS VDD 271 620 657 ICV_22 $T=117300 51680 1 0 $X=117110 $Y=48720
X1176 VSS VDD 301 510 301 ICV_22 $T=123280 62560 1 0 $X=123090 $Y=59600
X1177 VSS VDD 625 672 704 ICV_22 $T=125120 127840 1 0 $X=124930 $Y=124880
X1178 VSS VDD 617 677 617 ICV_22 $T=126500 127840 0 0 $X=126310 $Y=127600
X1179 VSS VDD 286 558 760 ICV_22 $T=133400 138720 1 0 $X=133210 $Y=135760
X1180 VSS VDD 387 289 387 ICV_22 $T=140300 73440 0 0 $X=140110 $Y=73200
X1181 VSS VDD PAR_IN4<12> 88 81 80 PAR_IN4<12> ICV_23 $T=7820 144160 0 0 $X=7630 $Y=143920
X1182 VSS VDD PAR_IN3<1> 101 85 91 PAR_IN3<1> ICV_23 $T=9660 116960 0 0 $X=9470 $Y=116720
X1183 VSS VDD PAR_IN8<7> 147 138 137 PAR_IN8<7> ICV_23 $T=19780 111520 0 0 $X=19590 $Y=111280
X1184 VSS VDD PAR_IN7<4> 230 244 164 PAR_IN7<4> ICV_23 $T=41400 149600 0 0 $X=41210 $Y=149360
X1185 VSS VDD PAR_IN8<4> 235 112 207 PAR_IN8<4> ICV_23 $T=46460 29920 0 0 $X=46270 $Y=29680
X1186 VSS VDD 342 344 342 336 PAR_IN2<9> ICV_23 $T=61180 138720 1 0 $X=60990 $Y=135760
X1187 VSS VDD COUNT<2> 361 319 353 407 ICV_23 $T=67160 106080 0 0 $X=66970 $Y=105840
X1188 VSS VDD PAR_IN8<6> 459 465 348 PAR_IN8<6> ICV_23 $T=77740 73440 0 0 $X=77550 $Y=73200
X1189 VSS VDD 228 528 457 228 PAR_IN3<22> ICV_23 $T=89240 106080 1 0 $X=89050 $Y=103120
X1190 VSS VDD 537 423 556 228 PAR_IN3<6> ICV_23 $T=92920 95200 1 0 $X=92730 $Y=92240
X1191 VSS VDD PAR_IN8<15> 580 148 432 PAR_IN8<15> ICV_23 $T=97980 122400 0 0 $X=97790 $Y=122160
X1192 VSS VDD 91 508 627 432 PAR_IN8<24> ICV_23 $T=105340 133280 1 0 $X=105150 $Y=130320
X1193 VSS VDD 647 636 647 654 PAR_IN2<10> ICV_23 $T=116840 111520 1 0 $X=116650 $Y=108560
X1194 VSS VDD 670 529 670 677 PAR_IN7<1> ICV_23 $T=117760 122400 1 0 $X=117570 $Y=119440
X1195 VSS VDD PAR_IN8<27> 732 695 137 PAR_IN8<27> ICV_23 $T=126040 29920 0 0 $X=125850 $Y=29680
X1196 VSS VDD PAR_IN2<30> 706 725 395 PAR_IN2<30> ICV_23 $T=126040 84320 0 0 $X=125850 $Y=84080
X1197 VSS VDD PAR_IN2<2> 729 738 654 PAR_IN2<2> ICV_23 $T=134780 95200 0 0 $X=134590 $Y=94960
X1198 VSS VDD 732 780 767 513 PAR_IN7<27> ICV_23 $T=135240 35360 1 0 $X=135050 $Y=32400
X1199 VSS VDD 667 753 667 653 PAR_IN4<23> ICV_23 $T=135240 100640 1 0 $X=135050 $Y=97680
X1200 VSS VDD PAR_IN4<23> 518 795 145 PAR_IN8<5> ICV_23 $T=138460 95200 1 0 $X=138270 $Y=92240
X1201 VSS VDD 395 752 774 387 PAR_IN3<28> ICV_23 $T=138920 133280 1 0 $X=138730 $Y=130320
X1202 VSS VDD 69 130 146 ICV_24 $T=35880 51680 1 0 $X=35690 $Y=48720
X1203 VSS VDD 243 257 229 ICV_24 $T=44620 122400 0 0 $X=44430 $Y=122160
X1204 VSS VDD PAR_IN3<13> 293 298 ICV_24 $T=52900 19040 0 0 $X=52710 $Y=18800
X1205 VSS VDD COUNT<2> 312 313 ICV_24 $T=54740 111520 0 0 $X=54550 $Y=111280
X1206 VSS VDD 319 407 353 ICV_24 $T=69000 106080 1 0 $X=68810 $Y=103120
X1207 VSS VDD 469 523 525 ICV_24 $T=91080 29920 0 0 $X=90890 $Y=29680
X1208 VSS VDD 227 59 512 ICV_24 $T=91080 106080 0 0 $X=90890 $Y=105840
X1209 VSS VDD 572 588 590 ICV_24 $T=100740 51680 0 0 $X=100550 $Y=51440
X1210 VSS VDD 609 405 636 ICV_24 $T=106260 95200 1 0 $X=106070 $Y=92240
X1211 VSS VDD 763 513 772 ICV_24 $T=135240 29920 1 0 $X=135050 $Y=26960
X1212 VSS VDD 285 745 381 ICV_24 $T=136620 57120 0 0 $X=136430 $Y=56880
X1213 VSS VDD 774 PAR_IN3<28> 387 ICV_24 $T=138920 127840 0 0 $X=138730 $Y=127600
X1214 VSS VDD PAR_IN2<1> 66 85 PAR_IN2<1> ICV_25 $T=8280 122400 0 0 $X=8090 $Y=122160
X1215 VSS VDD 83 161 177 83 ICV_25 $T=24380 24480 0 0 $X=24190 $Y=24240
X1216 VSS VDD 69 133 7 184 ICV_25 $T=26680 51680 0 0 $X=26490 $Y=51440
X1217 VSS VDD PAR_IN6<21> 59 280 PAR_IN6<21> ICV_25 $T=49220 100640 0 0 $X=49030 $Y=100400
X1218 VSS VDD COUNT<0> 37 232 COUNT<0> ICV_25 $T=50140 73440 0 0 $X=49950 $Y=73200
X1219 VSS VDD PAR_IN2<31> 290 315 PAR_IN2<31> ICV_25 $T=54740 13600 0 0 $X=54550 $Y=13360
X1220 VSS VDD PAR_IN5<17> 127 390 PAR_IN5<17> ICV_25 $T=65780 40800 0 0 $X=65590 $Y=40560
X1221 VSS VDD PAR_IN8<22> 373 480 PAR_IN8<22> ICV_25 $T=80960 106080 0 0 $X=80770 $Y=105840
X1222 VSS VDD PAR_IN5<14> 271 466 PAR_IN5<14> ICV_25 $T=82800 57120 0 0 $X=82610 $Y=56880
X1223 VSS VDD PAR_IN2<13> 336 298 PAR_IN2<13> ICV_25 $T=91080 19040 0 0 $X=90890 $Y=18800
X1224 VSS VDD PAR_IN7<15> 558 545 80 ICV_25 $T=97060 133280 1 0 $X=96870 $Y=130320
X1225 VSS VDD PAR_IN5<3> 563 553 513 ICV_25 $T=97060 155040 1 0 $X=96870 $Y=152080
X1226 VSS VDD PAR_IN6<22> 625 624 PAR_IN6<22> ICV_25 $T=110860 35360 0 0 $X=110670 $Y=35120
X1227 VSS VDD PAR_IN5<0> 67 648 PAR_IN5<0> ICV_25 $T=110860 149600 0 0 $X=110670 $Y=149360
X1228 VSS VDD PAR_IN5<27> 563 695 PAR_IN7<30> ICV_25 $T=119140 29920 0 0 $X=118950 $Y=29680
X1229 VSS VDD PAR_IN6<11> 437 766 796 ICV_25 $T=138000 78880 1 0 $X=137810 $Y=75920
X1230 VSS VDD PAR_IN7<9> 617 342 PAR_IN7<9> ICV_25 $T=138460 138720 0 0 $X=138270 $Y=138480
X1231 VSS VDD PAR_IN4<14> 754 559 PAR_IN4<14> ICV_25 $T=138920 51680 0 0 $X=138730 $Y=51440
X1232 VSS VDD PAR_IN5<5> 89 795 PAR_IN5<5> ICV_25 $T=138920 89760 0 0 $X=138730 $Y=89520
X1233 VSS VDD 49 29 ICV_26 $T=6900 68000 1 0 $X=6710 $Y=65040
X1234 VSS VDD RESET 167 ICV_26 $T=25300 106080 0 0 $X=25110 $Y=105840
X1235 VSS VDD PAR_IN8<25> 207 ICV_26 $T=31740 155040 1 0 $X=31550 $Y=152080
X1236 VSS VDD 59 25 ICV_26 $T=43240 100640 0 0 $X=43050 $Y=100400
X1237 VSS VDD 303 PAR_IN1<14> ICV_26 $T=62100 51680 0 0 $X=61910 $Y=51440
X1238 VSS VDD 287 135 ICV_26 $T=62100 73440 0 0 $X=61910 $Y=73200
X1239 VSS VDD 395 366 ICV_26 $T=65780 116960 1 0 $X=65590 $Y=114000
X1240 VSS VDD 147 449 ICV_26 $T=76360 100640 1 0 $X=76170 $Y=97680
X1241 VSS VDD 341 481 ICV_26 $T=80500 111520 1 0 $X=80310 $Y=108560
X1242 VSS VDD COUNT<2> 488 ICV_26 $T=80960 68000 0 0 $X=80770 $Y=67760
X1243 VSS VDD 396 526 ICV_26 $T=89240 40800 1 0 $X=89050 $Y=37840
X1244 VSS VDD 493 PAR_IN4<17> ICV_26 $T=100740 46240 0 0 $X=100550 $Y=46000
X1245 VSS VDD PAR_IN5<6> 604 ICV_26 $T=103500 62560 0 0 $X=103310 $Y=62320
X1246 VSS VDD 722 286 ICV_26 $T=125120 138720 1 0 $X=124930 $Y=135760
X1247 VSS VDD 395 387 ICV_26 $T=132480 116960 1 0 $X=132290 $Y=114000
X1248 VSS VDD PAR_IN8<28> 207 ICV_26 $T=138920 78880 0 0 $X=138730 $Y=78640
X1249 VSS VDD 145 146 97 ICV_27 $T=22540 73440 0 0 $X=22350 $Y=73200
X1250 VSS VDD 29 69 100 ICV_27 $T=26220 62560 1 0 $X=26030 $Y=59600
X1251 VSS VDD 240 240 143 ICV_27 $T=42780 35360 0 0 $X=42590 $Y=35120
X1252 VSS VDD 293 282 258 ICV_27 $T=53360 78880 0 0 $X=53170 $Y=78640
X1253 VSS VDD 20 178 293 ICV_27 $T=53820 89760 1 0 $X=53630 $Y=86800
X1254 VSS VDD 356 340 374 ICV_27 $T=63940 62560 1 0 $X=63750 $Y=59600
X1255 VSS VDD 282 282 66 ICV_27 $T=100280 62560 0 0 $X=100090 $Y=62320
X1256 VSS VDD 627 602 181 ICV_27 $T=110400 127840 1 0 $X=110210 $Y=124880
X1257 VSS VDD 604 374 457 ICV_27 $T=121440 73440 0 0 $X=121250 $Y=73200
X1258 VSS VDD 558 558 513 ICV_27 $T=138460 144160 1 0 $X=138270 $Y=141200
X1259 VSS VDD 161 165 ICV_28 $T=26220 29920 1 0 $X=26030 $Y=26960
X1260 VSS VDD PAR_IN1<10> 163 ICV_28 $T=39100 122400 0 0 $X=38910 $Y=122160
X1261 VSS VDD SAMPLE_COUNT<3> 234 ICV_28 $T=40020 73440 1 0 $X=39830 $Y=70480
X1262 VSS VDD 178 249 ICV_28 $T=42320 144160 1 0 $X=42130 $Y=141200
X1263 VSS VDD 215 268 ICV_28 $T=49220 62560 1 0 $X=49030 $Y=59600
X1264 VSS VDD PAR_IN3<31> 315 ICV_28 $T=57040 13600 1 0 $X=56850 $Y=10640
X1265 VSS VDD PAR_IN2<11> 272 ICV_28 $T=66240 13600 0 0 $X=66050 $Y=13360
X1266 VSS VDD PAR_IN2<21> 293 ICV_28 $T=82340 19040 0 0 $X=82150 $Y=18800
X1267 VSS VDD PAR_IN1<0> 383 ICV_28 $T=83720 144160 0 0 $X=83530 $Y=143920
X1268 VSS VDD PAR_IN4<21> 468 ICV_28 $T=97980 24480 1 0 $X=97790 $Y=21520
X1269 VSS VDD 66 528 ICV_28 $T=97980 111520 1 0 $X=97790 $Y=108560
X1270 VSS VDD 544 580 ICV_28 $T=106260 122400 0 0 $X=106070 $Y=122160
X1271 VSS VDD PAR_IN8<24> 432 ICV_28 $T=109940 127840 0 0 $X=109750 $Y=127600
X1272 VSS VDD PAR_IN1<21> 264 ICV_28 $T=110400 29920 0 0 $X=110210 $Y=29680
X1273 VSS VDD PAR_IN7<31> 715 ICV_28 $T=126500 24480 1 0 $X=126310 $Y=21520
X1274 VSS VDD 653 667 ICV_28 $T=136620 106080 1 0 $X=136430 $Y=103120
X1275 VSS VDD PAR_IN6<0> 762 ICV_28 $T=137540 19040 0 0 $X=137350 $Y=18800
X1276 VSS VDD 4 56 64 76 ICV_29 $T=10120 46240 1 0 $X=9930 $Y=43280
X1277 VSS VDD PAR_IN7<8> PAR_IN5<8> 140 188 ICV_29 $T=23920 138720 0 0 $X=23730 $Y=138480
X1278 VSS VDD 290 PAR_IN2<7> 290 316 ICV_29 $T=52900 24480 0 0 $X=52710 $Y=24240
X1279 VSS VDD 437 PAR_IN6<5> 437 575 ICV_29 $T=95680 155040 0 0 $X=95490 $Y=154800
X1280 VSS VDD 563 PAR_IN5<11> 563 626 ICV_29 $T=104880 73440 0 0 $X=104690 $Y=73200
X1281 VSS VDD 301 PAR_IN3<10> 301 635 ICV_29 $T=105800 89760 0 0 $X=105610 $Y=89520
X1282 VSS VDD 343 PAR_IN4<10> 343 647 ICV_29 $T=108560 116960 0 0 $X=108370 $Y=116720
X1283 VSS VDD 290 PAR_IN2<19> 290 693 ICV_29 $T=125120 89760 0 0 $X=124930 $Y=89520
X1284 VSS VDD PAR_IN6<30> PAR_IN6<30> 625 708 ICV_29 $T=127420 35360 0 0 $X=127230 $Y=35120
X1285 VSS VDD PAR_IN5<18> PAR_IN6<0> 546 768 ICV_29 $T=131560 19040 0 0 $X=131370 $Y=18800
X1286 VSS VDD 672 PAR_IN6<24> 672 734 ICV_29 $T=136160 122400 0 0 $X=135970 $Y=122160
X1287 VSS VDD PAR_IN3<0> PAR_IN2<0> 395 788 ICV_29 $T=137080 133280 0 0 $X=136890 $Y=133040
X1288 VSS VDD 121 88 94 128 VDD 163 VSS sky130_fd_sc_hd__or4_4 $T=21160 133280 1 0 $X=20970 $Y=130320
X1289 VSS VDD 182 175 187 156 VDD 196 VSS sky130_fd_sc_hd__or4_4 $T=28060 138720 1 0 $X=27870 $Y=135760
X1290 VSS VDD 173 93 208 168 VDD 214 VSS sky130_fd_sc_hd__or4_4 $T=33120 149600 1 0 $X=32930 $Y=146640
X1291 VSS VDD 223 COMPLETE COUNT<5> SAMPLE_COUNT<3> VDD 234 VSS sky130_fd_sc_hd__or4_4 $T=38640 73440 0 0 $X=38450 $Y=73200
X1292 VSS VDD 230 92 235 238 VDD 245 VSS sky130_fd_sc_hd__or4_4 $T=40480 138720 0 0 $X=40290 $Y=138480
X1293 VSS VDD 180 256 70 261 VDD 287 VSS sky130_fd_sc_hd__or4_4 $T=49680 78880 1 0 $X=49490 $Y=75920
X1294 VSS VDD 344 294 354 324 VDD 323 VSS sky130_fd_sc_hd__or4_4 $T=62560 149600 1 0 $X=62370 $Y=146640
X1295 VSS VDD 226 359 347 363 VDD 377 VSS sky130_fd_sc_hd__or4_4 $T=63940 29920 1 0 $X=63750 $Y=26960
X1296 VSS VDD 71 414 404 426 VDD 458 VSS sky130_fd_sc_hd__or4_4 $T=77280 40800 1 0 $X=77090 $Y=37840
X1297 VSS VDD 449 454 147 346 VDD 447 VSS sky130_fd_sc_hd__or4_4 $T=78660 100640 0 0 $X=78470 $Y=100400
X1298 VSS VDD 386 446 462 429 VDD 400 VSS sky130_fd_sc_hd__or4_4 $T=80040 57120 1 0 $X=79850 $Y=54160
X1299 VSS VDD 352 423 459 430 VDD 407 VSS sky130_fd_sc_hd__or4_4 $T=80040 95200 0 0 $X=79850 $Y=94960
X1300 VSS VDD 494 522 169 442 VDD 525 VSS sky130_fd_sc_hd__or4_4 $T=91080 24480 0 0 $X=90890 $Y=24240
X1301 VSS VDD 524 502 529 101 VDD 512 VSS sky130_fd_sc_hd__or4_4 $T=92000 116960 0 0 $X=91810 $Y=116720
X1302 VSS VDD 508 507 538 388 VDD 335 VSS sky130_fd_sc_hd__or4_4 $T=92000 138720 1 0 $X=91810 $Y=135760
X1303 VSS VDD 518 516 547 288 VDD 536 VSS sky130_fd_sc_hd__or4_4 $T=94760 84320 1 0 $X=94570 $Y=81360
X1304 VSS VDD 570 528 571 567 VDD 450 VSS sky130_fd_sc_hd__or4_4 $T=99360 106080 0 0 $X=99170 $Y=105840
X1305 VSS VDD 578 587 445 579 VDD 509 VSS sky130_fd_sc_hd__or4_4 $T=105340 40800 1 0 $X=105150 $Y=37840
X1306 VSS VDD 572 595 588 590 VDD 550 VSS sky130_fd_sc_hd__or4_4 $T=105340 57120 1 0 $X=105150 $Y=54160
X1307 VSS VDD 586 585 582 399 VDD 517 VSS sky130_fd_sc_hd__or4_4 $T=105340 73440 1 0 $X=105150 $Y=70480
X1308 VSS VDD 574 591 580 544 VDD 530 VSS sky130_fd_sc_hd__or4_4 $T=105340 127840 1 0 $X=105150 $Y=124880
X1309 VSS VDD 631 640 630 321 VDD 474 VSS sky130_fd_sc_hd__or4_4 $T=109940 24480 0 0 $X=109750 $Y=24240
X1310 VSS VDD 609 405 610 636 VDD 274 VSS sky130_fd_sc_hd__or4_4 $T=109940 95200 0 0 $X=109750 $Y=94960
X1311 VSS VDD 634 637 292 622 VDD 237 VSS sky130_fd_sc_hd__or4_4 $T=109940 106080 0 0 $X=109750 $Y=105840
X1312 VSS VDD 655 650 633 659 VDD 534 VSS sky130_fd_sc_hd__or4_4 $T=115460 73440 1 0 $X=115270 $Y=70480
X1313 VSS VDD 706 674 705 696 VDD 416 VSS sky130_fd_sc_hd__or4_4 $T=124200 51680 1 0 $X=124010 $Y=48720
X1314 VSS VDD 707 727 698 726 VDD 471 VSS sky130_fd_sc_hd__or4_4 $T=127880 111520 0 0 $X=127690 $Y=111280
X1315 VSS VDD 731 710 730 720 VDD 357 VSS sky130_fd_sc_hd__or4_4 $T=128800 62560 0 0 $X=128610 $Y=62320
X1316 VSS VDD 729 728 381 745 VDD 320 VSS sky130_fd_sc_hd__or4_4 $T=131560 57120 0 0 $X=131370 $Y=56880
X1317 VSS VDD 683 753 742 746 VDD 492 VSS sky130_fd_sc_hd__or4_4 $T=133400 95200 1 0 $X=133210 $Y=92240
X1318 VSS VDD 747 736 628 752 VDD 477 VSS sky130_fd_sc_hd__or4_4 $T=133400 127840 1 0 $X=133210 $Y=124880
X1319 VSS VDD 687 722 714 760 VDD 453 VSS sky130_fd_sc_hd__or4_4 $T=133400 144160 1 0 $X=133210 $Y=141200
X1320 VSS VDD 732 763 780 772 VDD 549 VSS sky130_fd_sc_hd__or4_4 $T=137080 29920 0 0 $X=136890 $Y=29680
X1321 VSS VDD PAR_IN4<8> 181 ICV_30 $T=23460 122400 0 0 $X=23270 $Y=122160
X1322 VSS VDD RESET 177 ICV_30 $T=23920 19040 0 0 $X=23730 $Y=18800
X1323 VSS VDD 320 326 ICV_30 $T=56120 73440 1 0 $X=55930 $Y=70480
X1324 VSS VDD 382 COUNT<4> ICV_30 $T=65780 122400 0 0 $X=65590 $Y=122160
X1325 VSS VDD 383 PAR_IN1<25> ICV_30 $T=74520 144160 0 0 $X=74330 $Y=143920
X1326 VSS VDD 491 202 ICV_30 $T=84640 62560 0 0 $X=84450 $Y=62320
X1327 VSS VDD 654 PAR_IN2<26> ICV_30 $T=112700 111520 0 0 $X=112510 $Y=111280
X1328 VSS VDD 648 437 ICV_30 $T=114080 155040 1 0 $X=113890 $Y=152080
X1329 VSS VDD 710 720 ICV_30 $T=123740 62560 0 0 $X=123550 $Y=62320
X1330 VSS VDD 738 654 ICV_30 $T=129720 95200 0 0 $X=129530 $Y=94960
X1331 VSS VDD PAR_IN6<23> 643 ICV_30 $T=136620 149600 0 0 $X=136430 $Y=149360
X1332 VSS VDD 69 ICV_31 $T=6900 62560 1 0 $X=6710 $Y=59600
X1333 VSS VDD PAR_IN4<25> ICV_31 $T=6900 149600 0 0 $X=6710 $Y=149360
X1334 VSS VDD RESET ICV_31 $T=11040 106080 0 0 $X=10850 $Y=105840
X1335 VSS VDD 64 ICV_31 $T=16100 62560 1 0 $X=15910 $Y=59600
X1336 VSS VDD 118 ICV_31 $T=16100 84320 1 0 $X=15910 $Y=81360
X1337 VSS VDD PAR_IN5<15> ICV_31 $T=16560 122400 0 0 $X=16370 $Y=122160
X1338 VSS VDD 89 ICV_31 $T=18400 29920 0 0 $X=18210 $Y=29680
X1339 VSS VDD 100 ICV_31 $T=18400 62560 0 0 $X=18210 $Y=62320
X1340 VSS VDD 133 ICV_31 $T=23000 51680 0 0 $X=22810 $Y=51440
X1341 VSS VDD 184 ICV_31 $T=29900 46240 0 0 $X=29710 $Y=46000
X1342 VSS VDD 194 ICV_31 $T=31280 73440 1 0 $X=31090 $Y=70480
X1343 VSS VDD 165 ICV_31 $T=31280 100640 1 0 $X=31090 $Y=97680
X1344 VSS VDD 93 ICV_31 $T=31280 144160 1 0 $X=31090 $Y=141200
X1345 VSS VDD 133 ICV_31 $T=32200 57120 1 0 $X=32010 $Y=54160
X1346 VSS VDD 207 ICV_31 $T=32200 138720 1 0 $X=32010 $Y=135760
X1347 VSS VDD 115 ICV_31 $T=34040 57120 0 0 $X=33850 $Y=56880
X1348 VSS VDD COUNT<3> ICV_31 $T=37260 116960 0 0 $X=37070 $Y=116720
X1349 VSS VDD 143 ICV_31 $T=44160 46240 1 0 $X=43970 $Y=43280
X1350 VSS VDD 56 ICV_31 $T=44160 51680 1 0 $X=43970 $Y=48720
X1351 VSS VDD SAMPLE_COUNT<0> ICV_31 $T=46000 35360 0 0 $X=45810 $Y=35120
X1352 VSS VDD PAR_IN3<9> ICV_31 $T=48760 149600 0 0 $X=48570 $Y=149360
X1353 VSS VDD 258 ICV_31 $T=52900 68000 1 0 $X=52710 $Y=65040
X1354 VSS VDD 305 ICV_31 $T=54740 106080 1 0 $X=54550 $Y=103120
X1355 VSS VDD 309 ICV_31 $T=57040 133280 1 0 $X=56850 $Y=130320
X1356 VSS VDD COUNT<4> ICV_31 $T=57960 68000 0 0 $X=57770 $Y=67760
X1357 VSS VDD 214 ICV_31 $T=68080 144160 1 0 $X=67890 $Y=141200
X1358 VSS VDD 202 ICV_31 $T=74520 89760 0 0 $X=74330 $Y=89520
X1359 VSS VDD 346 ICV_31 $T=74980 100640 0 0 $X=74790 $Y=100400
X1360 VSS VDD 392 ICV_31 $T=78660 78880 0 0 $X=78470 $Y=78640
X1361 VSS VDD 469 ICV_31 $T=80500 35360 0 0 $X=80310 $Y=35120
X1362 VSS VDD 118 ICV_31 $T=86020 68000 0 0 $X=85830 $Y=67760
X1363 VSS VDD PAR_IN1<1> ICV_31 $T=86020 111520 0 0 $X=85830 $Y=111280
X1364 VSS VDD 227 ICV_31 $T=86020 127840 0 0 $X=85830 $Y=127600
X1365 VSS VDD PAR_IN2<22> ICV_31 $T=94300 111520 0 0 $X=94110 $Y=111280
X1366 VSS VDD 392 ICV_31 $T=97060 78880 0 0 $X=96870 $Y=78640
X1367 VSS VDD PAR_IN3<15> ICV_31 $T=99820 127840 0 0 $X=99630 $Y=127600
X1368 VSS VDD PAR_IN7<28> ICV_31 $T=104420 133280 0 0 $X=104230 $Y=133040
X1369 VSS VDD 625 ICV_31 $T=107180 35360 0 0 $X=106990 $Y=35120
X1370 VSS VDD 611 ICV_31 $T=110860 100640 1 0 $X=110670 $Y=97680
X1371 VSS VDD PAR_IN5<31> ICV_31 $T=114080 13600 0 0 $X=113890 $Y=13360
X1372 VSS VDD PAR_IN5<1> ICV_31 $T=114080 19040 0 0 $X=113890 $Y=18800
X1373 VSS VDD 654 ICV_31 $T=114080 106080 0 0 $X=113890 $Y=105840
X1374 VSS VDD PAR_IN3<18> ICV_31 $T=128340 68000 0 0 $X=128150 $Y=67760
X1375 VSS VDD PAR_IN7<27> ICV_31 $T=133400 29920 0 0 $X=133210 $Y=29680
X1376 VSS VDD 558 ICV_31 $T=134780 138720 0 0 $X=134590 $Y=138480
X1377 VSS VDD 155 116 118 146 202 ICV_32 $T=24380 84320 0 0 $X=24190 $Y=84080
X1378 VSS VDD 261 298 293 PAR_IN3<13> 226 ICV_32 $T=52440 24480 1 0 $X=52250 $Y=21520
X1379 VSS VDD 346 316 289 PAR_IN3<7> 293 ICV_32 $T=61640 24480 1 0 $X=61450 $Y=21520
X1380 VSS VDD 363 371 89 PAR_IN5<20> 396 ICV_32 $T=64400 29920 0 0 $X=64210 $Y=29680
X1381 VSS VDD 354 389 102 PAR_IN8<9> PAR_IN6<9> ICV_32 $T=66700 149600 0 0 $X=66510 $Y=149360
X1382 VSS VDD 399 398 293 PAR_IN3<11> PAR_IN3<21> ICV_32 $T=69000 19040 0 0 $X=68810 $Y=18800
X1383 VSS VDD 404 114 145 PAR_IN8<29> 396 ICV_32 $T=78200 40800 0 0 $X=78010 $Y=40560
X1384 VSS VDD 570 480 66 PAR_IN2<22> PAR_IN7<22> ICV_32 $T=97980 111520 0 0 $X=97790 $Y=111280
X1385 VSS VDD 714 768 558 PAR_IN7<0> PAR_IN5<24> ICV_32 $T=136620 144160 0 0 $X=136430 $Y=143920
X1386 VSS VDD COUNT<0> 154 116 14 97 ICV_33 $T=23920 89760 0 0 $X=23730 $Y=89520
X1387 VSS VDD 140 168 106 178 PAR_IN3<25> ICV_33 $T=23920 149600 1 0 $X=23730 $Y=146640
X1388 VSS VDD 146 180 150 145 PAR_IN8<13> ICV_33 $T=25760 78880 1 0 $X=25570 $Y=75920
X1389 VSS VDD PAR_IN1<4> 294 304 178 PAR_IN3<9> ICV_33 $T=52440 149600 0 0 $X=52250 $Y=149360
X1390 VSS VDD 558 502 493 181 PAR_IN4<1> ICV_33 $T=90620 127840 1 0 $X=90430 $Y=124880
X1391 VSS VDD 563 507 304 80 PAR_IN4<24> ICV_33 $T=91080 149600 1 0 $X=90890 $Y=146640
X1392 VSS VDD 457 359 493 59 PAR_IN6<20> ICV_33 $T=92460 100640 0 0 $X=92270 $Y=100400
X1393 VSS VDD 560 544 537 59 PAR_IN6<15> ICV_33 $T=94300 100640 1 0 $X=94110 $Y=97680
X1394 VSS VDD 625 628 606 558 PAR_IN7<28> ICV_33 $T=108100 133280 0 0 $X=107910 $Y=133040
X1395 VSS VDD 705 674 457 510 PAR_IN3<30> ICV_33 $T=117760 46240 1 0 $X=117570 $Y=43280
X1396 VSS VDD 102 698 709 102 PAR_IN8<16> ICV_33 $T=122360 57120 0 0 $X=122170 $Y=56880
X1397 VSS VDD 625 705 708 617 PAR_IN7<30> ICV_33 $T=122820 35360 1 0 $X=122630 $Y=32400
X1398 VSS VDD 286 538 734 677 PAR_IN7<24> ICV_33 $T=127880 133280 0 0 $X=127690 $Y=133040
X1399 VSS VDD 510 710 374 510 PAR_IN3<18> ICV_33 $T=132020 68000 0 0 $X=131830 $Y=67760
X1400 VSS VDD 768 722 304 560 PAR_IN4<0> ICV_33 $T=134780 149600 1 0 $X=134590 $Y=146640
X1401 VSS VDD PAR_IN8<26> 726 338 387 PAR_IN3<16> ICV_33 $T=136160 111520 0 0 $X=135970 $Y=111280
X1402 VSS VDD 667 763 667 653 PAR_IN4<27> ICV_33 $T=136620 35360 0 0 $X=136430 $Y=35120
X1403 VSS VDD 78 ICV_34 $T=11500 84320 0 0 $X=11310 $Y=84080
X1404 VSS VDD 108 ICV_34 $T=14260 100640 1 0 $X=14070 $Y=97680
X1405 VSS VDD 79 ICV_34 $T=14260 111520 0 0 $X=14070 $Y=111280
X1406 VSS VDD 110 ICV_34 $T=14720 106080 1 0 $X=14530 $Y=103120
X1407 VSS VDD 49 ICV_34 $T=14720 111520 1 0 $X=14530 $Y=108560
X1408 VSS VDD 103 ICV_34 $T=15180 122400 1 0 $X=14990 $Y=119440
X1409 VSS VDD PAR_IN5<21> ICV_34 $T=28060 13600 0 0 $X=27870 $Y=13360
X1410 VSS VDD 197 ICV_34 $T=37720 155040 1 0 $X=37530 $Y=152080
X1411 VSS VDD 215 ICV_34 $T=40020 57120 0 0 $X=39830 $Y=56880
X1412 VSS VDD 223 ICV_34 $T=41400 78880 1 0 $X=41210 $Y=75920
X1413 VSS VDD 164 ICV_34 $T=43240 149600 1 0 $X=43050 $Y=146640
X1414 VSS VDD 244 ICV_34 $T=43240 155040 1 0 $X=43050 $Y=152080
X1415 VSS VDD 196 ICV_34 $T=43700 127840 0 0 $X=43510 $Y=127600
X1416 VSS VDD 337 ICV_34 $T=61640 78880 1 0 $X=61450 $Y=75920
X1417 VSS VDD 373 ICV_34 $T=69000 95200 1 0 $X=68810 $Y=92240
X1418 VSS VDD 403 ICV_34 $T=69000 100640 1 0 $X=68810 $Y=97680
X1419 VSS VDD 354 ICV_34 $T=69920 144160 0 0 $X=69730 $Y=143920
X1420 VSS VDD 319 ICV_34 $T=70840 122400 1 0 $X=70650 $Y=119440
X1421 VSS VDD 397 ICV_34 $T=71300 127840 0 0 $X=71110 $Y=127600
X1422 VSS VDD 359 ICV_34 $T=71760 24480 0 0 $X=71570 $Y=24240
X1423 VSS VDD 281 ICV_34 $T=78660 116960 0 0 $X=78470 $Y=116720
X1424 VSS VDD 431 ICV_34 $T=98440 19040 1 0 $X=98250 $Y=16080
X1425 VSS VDD 431 ICV_34 $T=98440 89760 1 0 $X=98250 $Y=86800
X1426 VSS VDD 516 ICV_34 $T=98900 78880 1 0 $X=98710 $Y=75920
X1427 VSS VDD 336 ICV_34 $T=98900 138720 1 0 $X=98710 $Y=135760
X1428 VSS VDD 413 ICV_34 $T=99820 13600 1 0 $X=99630 $Y=10640
X1429 VSS VDD PAR_IN5<11> ICV_34 $T=110860 73440 0 0 $X=110670 $Y=73200
X1430 VSS VDD PAR_IN2<17> ICV_34 $T=111320 51680 0 0 $X=111130 $Y=51440
X1431 VSS VDD 602 ICV_34 $T=112240 122400 0 0 $X=112050 $Y=122160
X1432 VSS VDD 635 ICV_34 $T=113160 89760 1 0 $X=112970 $Y=86800
X1433 VSS VDD 667 ICV_34 $T=117300 35360 1 0 $X=117110 $Y=32400
X1434 VSS VDD 563 ICV_34 $T=118220 29920 1 0 $X=118030 $Y=26960
X1435 VSS VDD 457 ICV_34 $T=127420 46240 1 0 $X=127230 $Y=43280
X1436 VSS VDD 67 ICV_34 $T=128340 13600 1 0 $X=128150 $Y=10640
X1437 VSS VDD 374 ICV_34 $T=135700 73440 1 0 $X=135510 $Y=70480
X1438 VSS 81 PAR_IN2<25> 80 66 ICV_35 $T=9660 149600 1 0 $X=9470 $Y=146640
X1439 VSS 83 97 76 49 ICV_35 $T=10580 29920 1 0 $X=10390 $Y=26960
X1440 VSS 121 128 94 88 ICV_35 $T=18400 127840 0 0 $X=18210 $Y=127600
X1441 VSS 170 4 157 198 ICV_35 $T=25760 35360 0 0 $X=25570 $Y=35120
X1442 VSS PAR_IN5<13> RESET 174 RESET ICV_35 $T=26220 29920 0 0 $X=26030 $Y=29680
X1443 VSS 158 187 175 182 ICV_35 $T=26220 133280 1 0 $X=26030 $Y=130320
X1444 VSS 168 208 173 PAR_IN3<4> ICV_35 $T=34960 144160 0 0 $X=34770 $Y=143920
X1445 VSS 215 130 130 211 ICV_35 $T=51520 46240 0 0 $X=51330 $Y=46000
X1446 VSS PAR_IN2<24> 258 324 PAR_IN1<6> ICV_35 $T=54280 144160 0 0 $X=54090 $Y=143920
X1447 VSS 89 371 363 347 ICV_35 $T=64400 24480 0 0 $X=64210 $Y=24240
X1448 VSS 21 25 401 23 ICV_35 $T=66700 78880 1 0 $X=66510 $Y=75920
X1449 VSS 446 373 466 462 ICV_35 $T=78200 51680 1 0 $X=78010 $Y=48720
X1450 VSS PAR_IN6<7> 437 486 PAR_IN7<7> ICV_35 $T=82340 149600 0 0 $X=82150 $Y=149360
X1451 VSS 474 490 458 509 ICV_35 $T=83720 35360 1 0 $X=83530 $Y=32400
X1452 VSS 186 101 432 548 ICV_35 $T=90160 116960 1 0 $X=89970 $Y=114000
X1453 VSS 578 587 579 445 ICV_35 $T=100740 35360 0 0 $X=100550 $Y=35120
X1454 VSS 582 399 137 PAR_IN8<19> ICV_35 $T=101200 68000 0 0 $X=101010 $Y=67760
X1455 VSS 667 PAR_IN3<19> 289 693 ICV_35 $T=116840 78880 1 0 $X=116650 $Y=75920
X1456 VSS 617 708 513 137 ICV_35 $T=122820 29920 1 0 $X=122630 $Y=26960
X1457 VSS PAR_IN4<6> 677 304 560 ICV_35 $T=125120 116960 0 0 $X=124930 $Y=116720
X1458 VSS 304 560 PAR_IN7<0> PAR_IN4<0> ICV_35 $T=129260 144160 0 0 $X=129070 $Y=143920
X1459 VSS PAR_IN2<19> 746 742 753 ICV_35 $T=131100 89760 0 0 $X=130910 $Y=89520
X1460 VSS 677 PAR_IN4<16> 560 304 ICV_35 $T=134320 106080 0 0 $X=134130 $Y=105840
X1461 VSS VDD ICV_36 $T=53360 35360 1 0 $X=53170 $Y=32400
X1462 VSS VDD ICV_36 $T=96140 40800 0 0 $X=95950 $Y=40560
X1463 VSS VDD ICV_36 $T=99820 116960 0 0 $X=99630 $Y=116720
X1464 VSS VDD ICV_36 $T=103960 84320 0 0 $X=103770 $Y=84080
X1465 VSS VDD ICV_36 $T=107180 40800 0 0 $X=106990 $Y=40560
X1466 VSS VDD ICV_36 $T=115000 62560 1 0 $X=114810 $Y=59600
X1467 VSS VDD ICV_36 $T=123280 78880 1 0 $X=123090 $Y=75920
X1468 VSS VDD ICV_36 $T=123280 149600 1 0 $X=123090 $Y=146640
X1469 VSS VDD ICV_37 $T=34040 155040 0 0 $X=33850 $Y=154800
X1470 VSS VDD ICV_37 $T=48300 155040 0 0 $X=48110 $Y=154800
X1471 VSS VDD ICV_37 $T=62560 13600 1 0 $X=62370 $Y=10640
X1472 VSS VDD ICV_37 $T=62560 155040 0 0 $X=62370 $Y=154800
X1473 VSS VDD ICV_37 $T=76820 155040 0 0 $X=76630 $Y=154800
X1474 VSS VDD ICV_37 $T=105340 155040 0 0 $X=105150 $Y=154800
X1475 VSS VDD ICV_37 $T=119600 155040 0 0 $X=119410 $Y=154800
X1476 VSS VDD ICV_37 $T=133860 13600 1 0 $X=133670 $Y=10640
X1477 VSS VDD ICV_37 $T=133860 155040 0 0 $X=133670 $Y=154800
X1478 VSS VDD 100 COUNT<1> ICV_38 $T=18400 100640 0 0 $X=18210 $Y=100400
X1479 VSS VDD 100 133 ICV_38 $T=20240 95200 0 0 $X=20050 $Y=94960
X1480 VSS VDD COUNT<1> 13 ICV_38 $T=26680 89760 1 0 $X=26490 $Y=86800
X1481 VSS VDD 227 224 ICV_38 $T=38180 127840 0 0 $X=37990 $Y=127600
X1482 VSS VDD PAR_IN1<18> 303 ICV_38 $T=52900 57120 0 0 $X=52710 $Y=56880
X1483 VSS VDD 332 336 ICV_38 $T=57960 29920 1 0 $X=57770 $Y=26960
X1484 VSS VDD 422 14 ICV_38 $T=72220 73440 0 0 $X=72030 $Y=73200
X1485 VSS VDD 518 535 ICV_38 $T=89240 84320 1 0 $X=89050 $Y=81360
X1486 VSS VDD 558 602 ICV_38 $T=112240 138720 0 0 $X=112050 $Y=138480
X1487 VSS VDD 140 PAR_IN8<30> ICV_38 $T=133400 84320 0 0 $X=133210 $Y=84080
X1488 VSS VDD 92 81 80 PAR_IN4<4> ICV_39 $T=10580 138720 1 0 $X=10390 $Y=135760
X1489 VSS VDD 169 176 145 PAR_IN8<21> ICV_39 $T=24380 19040 1 0 $X=24190 $Y=16080
X1490 VSS VDD 175 81 181 PAR_IN4<8> ICV_39 $T=24840 127840 1 0 $X=24650 $Y=124880
X1491 VSS VDD 226 231 181 PAR_IN4<20> ICV_39 $T=38640 19040 1 0 $X=38450 $Y=16080
X1492 VSS VDD 288 273 293 PAR_IN3<5> ICV_39 $T=51520 84320 1 0 $X=51330 $Y=81360
X1493 VSS VDD 321 315 289 PAR_IN3<31> ICV_39 $T=57040 19040 1 0 $X=56850 $Y=16080
X1494 VSS VDD 388 314 387 PAR_IN3<24> ICV_39 $T=66700 133280 0 0 $X=66510 $Y=133040
X1495 VSS VDD 386 366 395 PAR_IN2<14> ICV_39 $T=68080 111520 0 0 $X=67890 $Y=111280
X1496 VSS VDD 595 493 181 PAR_IN4<3> ICV_39 $T=108100 51680 1 0 $X=107910 $Y=48720
X1497 VSS VDD 582 626 137 PAR_IN8<11> ICV_39 $T=113620 68000 1 0 $X=113430 $Y=65040
X1498 VSS VDD 650 667 653 PAR_IN4<19> ICV_39 $T=117760 84320 1 0 $X=117570 $Y=81360
X1499 VSS VDD 683 652 145 PAR_IN8<23> ICV_39 $T=118680 89760 1 0 $X=118490 $Y=86800
X1500 VSS VDD 637 374 301 PAR_IN3<26> ICV_39 $T=122820 100640 0 0 $X=122630 $Y=100400
X1501 VSS VDD 707 699 677 PAR_IN7<16> ICV_39 $T=122820 106080 0 0 $X=122630 $Y=105840
X1502 VSS VDD 631 715 513 PAR_IN7<31> ICV_39 $T=126500 24480 0 0 $X=126310 $Y=24240
X1503 VSS VDD 720 762 620 PAR_IN5<18> ICV_39 $T=133400 24480 1 0 $X=133210 $Y=21520
X1504 VSS VDD 91 PAR_IN3<8> 156 141 91 PAR_IN3<8> ICV_40 $T=18860 144160 0 0 $X=18670 $Y=143920
X1505 VSS VDD 130 82 170 82 6 143 ICV_40 $T=20700 40800 0 0 $X=20510 $Y=40560
X1506 VSS VDD 111 PAR_IN7<25> 173 111 164 PAR_IN7<25> ICV_40 $T=20700 149600 0 0 $X=20510 $Y=149360
X1507 VSS VDD 141 PAR_IN3<25> 182 129 164 PAR_IN7<8> ICV_40 $T=22080 144160 1 0 $X=21890 $Y=141200
X1508 VSS VDD 260 PAR_IN7<26> 292 260 286 PAR_IN7<26> ICV_40 $T=48760 68000 0 0 $X=48570 $Y=67760
X1509 VSS VDD 319 PAR_IN8<10> 405 374 373 PAR_IN8<10> ICV_40 $T=65320 89760 0 0 $X=65130 $Y=89520
X1510 VSS VDD 429 PAR_IN8<14> 462 466 373 PAR_IN8<14> ICV_40 $T=76360 51680 0 0 $X=76170 $Y=51440
X1511 VSS VDD 431 PAR_IN4<29> 414 468 431 PAR_IN4<29> ICV_40 $T=76820 24480 0 0 $X=76630 $Y=24240
X1512 VSS VDD 396 455 494 280 77 PAR_IN7<21> ICV_40 $T=81880 29920 1 0 $X=81690 $Y=26960
X1513 VSS VDD 545 PAR_IN2<15> 574 545 336 PAR_IN2<15> ICV_40 $T=95220 133280 0 0 $X=95030 $Y=133040
X1514 VSS VDD 553 PAR_IN8<3> 572 553 137 PAR_IN8<3> ICV_40 $T=96140 144160 0 0 $X=95950 $Y=143920
X1515 VSS VDD 556 PAR_IN5<22> 567 621 620 PAR_IN5<22> ICV_40 $T=103960 100640 0 0 $X=103770 $Y=100400
X1516 VSS VDD 593 PAR_IN8<31> 630 629 432 PAR_IN8<31> ICV_40 $T=104880 19040 0 0 $X=104690 $Y=18800
X1517 VSS VDD 633 PAR_IN7<19> 655 688 77 PAR_IN7<19> ICV_40 $T=119140 68000 0 0 $X=118950 $Y=67760
X1518 VSS VDD 714 PAR_IN7<18> 730 701 286 PAR_IN7<18> ICV_40 $T=125580 138720 0 0 $X=125390 $Y=138480
X1519 VSS VDD 740 PAR_IN3<27> 696 776 620 PAR_IN5<30> ICV_40 $T=132020 40800 0 0 $X=131830 $Y=40560
X1520 VSS VDD 560 PAR_IN4<7> 454 667 653 PAR_IN4<7> ICV_40 $T=132940 100640 0 0 $X=132750 $Y=100400
X1521 VSS VDD 72 ICV_41 $T=6900 46240 0 0 $X=6710 $Y=46000
X1522 VSS VDD 26 ICV_41 $T=6900 62560 0 0 $X=6710 $Y=62320
X1523 VSS VDD 83 ICV_41 $T=11960 68000 1 0 $X=11770 $Y=65040
X1524 VSS VDD 166 ICV_41 $T=22540 78880 0 0 $X=22350 $Y=78640
X1525 VSS VDD 135 ICV_41 $T=29440 73440 0 0 $X=29250 $Y=73200
X1526 VSS VDD 247 ICV_41 $T=41860 95200 1 0 $X=41670 $Y=92240
X1527 VSS VDD 253 ICV_41 $T=43700 127840 1 0 $X=43510 $Y=124880
X1528 VSS VDD 289 ICV_41 $T=50600 13600 0 0 $X=50410 $Y=13360
X1529 VSS VDD PAR_IN2<20> ICV_41 $T=57500 29920 0 0 $X=57310 $Y=29680
X1530 VSS VDD 335 ICV_41 $T=57500 122400 0 0 $X=57310 $Y=122160
X1531 VSS VDD PAR_IN8<2> ICV_41 $T=62100 46240 0 0 $X=61910 $Y=46000
X1532 VSS VDD 22 ICV_41 $T=64860 84320 1 0 $X=64670 $Y=81360
X1533 VSS VDD PAR_IN8<29> ICV_41 $T=74060 40800 0 0 $X=73870 $Y=40560
X1534 VSS VDD PAR_IN1<23> ICV_41 $T=74520 106080 0 0 $X=74330 $Y=105840
X1535 VSS VDD PAR_IN1<30> ICV_41 $T=85560 51680 0 0 $X=85370 $Y=51440
X1536 VSS VDD 510 ICV_41 $T=86940 46240 1 0 $X=86750 $Y=43280
X1537 VSS VDD 137 ICV_41 $T=97520 144160 1 0 $X=97330 $Y=141200
X1538 VSS VDD PAR_IN6<12> ICV_41 $T=105340 144160 0 0 $X=105150 $Y=143920
X1539 VSS VDD PAR_IN6<17> ICV_41 $T=106720 13600 0 0 $X=106530 $Y=13360
X1540 VSS VDD PAR_IN5<26> ICV_41 $T=113160 100640 0 0 $X=112970 $Y=100400
X1541 VSS VDD 102 ICV_41 $T=115920 149600 1 0 $X=115730 $Y=146640
X1542 VSS VDD PAR_IN8<16> ICV_41 $T=118220 57120 0 0 $X=118030 $Y=56880
X1543 VSS VDD PAR_IN7<11> ICV_41 $T=129260 78880 0 0 $X=129070 $Y=78640
X1544 VSS VDD PAR_IN3<16> ICV_41 $T=132020 111520 0 0 $X=131830 $Y=111280
X1545 VSS VDD PAR_IN4<27> ICV_41 $T=132480 35360 0 0 $X=132290 $Y=35120
X1546 VSS VDD ICV_42 $T=19780 144160 1 0 $X=19590 $Y=141200
X1547 VSS VDD ICV_42 $T=33580 13600 0 0 $X=33390 $Y=13360
X1548 VSS VDD ICV_42 $T=33580 116960 0 0 $X=33390 $Y=116720
X1549 VSS VDD ICV_42 $T=33580 133280 0 0 $X=33390 $Y=133040
X1550 VSS VDD ICV_42 $T=61640 24480 0 0 $X=61450 $Y=24240
X1551 VSS VDD ICV_42 $T=61640 29920 0 0 $X=61450 $Y=29680
X1552 VSS VDD ICV_42 $T=61640 62560 0 0 $X=61450 $Y=62320
X1553 VSS VDD ICV_42 $T=61640 111520 0 0 $X=61450 $Y=111280
X1554 VSS VDD ICV_42 $T=75900 46240 1 0 $X=75710 $Y=43280
X1555 VSS VDD ICV_42 $T=75900 51680 1 0 $X=75710 $Y=48720
X1556 VSS VDD ICV_42 $T=89700 13600 0 0 $X=89510 $Y=13360
X1557 VSS VDD ICV_42 $T=89700 62560 0 0 $X=89510 $Y=62320
X1558 VSS VDD ICV_42 $T=89700 100640 0 0 $X=89510 $Y=100400
X1559 VSS VDD ICV_42 $T=89700 116960 0 0 $X=89510 $Y=116720
X1560 VSS VDD ICV_42 $T=89700 133280 0 0 $X=89510 $Y=133040
X1561 VSS VDD ICV_42 $T=103960 95200 1 0 $X=103770 $Y=92240
X1562 VSS VDD ICV_42 $T=103960 111520 1 0 $X=103770 $Y=108560
X1563 VSS VDD ICV_42 $T=132020 62560 1 0 $X=131830 $Y=59600
X1564 VSS VDD ICV_42 $T=132020 106080 1 0 $X=131830 $Y=103120
X1565 VSS VDD ICV_42 $T=132020 149600 1 0 $X=131830 $Y=146640
X1566 VSS 6 82 ICV_43 $T=19780 46240 1 0 $X=19590 $Y=43280
X1567 VSS 7 6 ICV_43 $T=19780 51680 1 0 $X=19590 $Y=48720
X1568 VSS COUNT<5> COMPLETE ICV_43 $T=33580 73440 0 0 $X=33390 $Y=73200
X1569 VSS 14 11 ICV_43 $T=33580 95200 0 0 $X=33390 $Y=94960
X1570 VSS RESET 171 ICV_43 $T=33580 100640 0 0 $X=33390 $Y=100400
X1571 VSS 259 278 ICV_43 $T=47840 111520 1 0 $X=47650 $Y=108560
X1572 VSS 262 242 ICV_43 $T=47840 116960 1 0 $X=47650 $Y=114000
X1573 VSS 319 24 ICV_43 $T=61640 78880 0 0 $X=61450 $Y=78640
X1574 VSS 341 308 ICV_43 $T=61640 122400 0 0 $X=61450 $Y=122160
X1575 VSS 344 PAR_IN8<9> ICV_43 $T=61640 149600 0 0 $X=61450 $Y=149360
X1576 VSS 227 410 ICV_43 $T=75900 89760 1 0 $X=75710 $Y=86800
X1577 VSS 401 454 ICV_43 $T=75900 106080 1 0 $X=75710 $Y=103120
X1578 VSS 437 441 ICV_43 $T=75900 155040 1 0 $X=75710 $Y=152080
X1579 VSS PAR_IN4<1> 493 ICV_43 $T=89700 122400 0 0 $X=89510 $Y=122160
X1580 VSS 413 401 ICV_43 $T=91080 13600 1 0 $X=90890 $Y=10640
X1581 VSS PAR_IN4<11> 431 ICV_43 $T=103960 78880 1 0 $X=103770 $Y=75920
X1582 VSS 591 574 ICV_43 $T=103960 122400 1 0 $X=103770 $Y=119440
X1583 VSS PAR_IN4<31> 653 ICV_43 $T=117760 35360 0 0 $X=117570 $Y=35120
X1584 VSS PAR_IN8<23> 145 ICV_43 $T=117760 84320 0 0 $X=117570 $Y=84080
X1585 VSS PAR_IN2<10> PAR_IN7<16> ICV_43 $T=117760 106080 0 0 $X=117570 $Y=105840
X1586 VSS 77 766 ICV_43 $T=132020 84320 1 0 $X=131830 $Y=81360
X1587 VSS 683 89 ICV_43 $T=132020 89760 1 0 $X=131830 $Y=86800
X1588 VSS VDD SAMPLE_COUNT<3> 146 ICV_44 $T=33580 68000 0 0 $X=33390 $Y=67760
X1589 VSS VDD 102 137 ICV_44 $T=33580 138720 0 0 $X=33390 $Y=138480
X1590 VSS VDD SAMPLE_COUNT<1> 211 ICV_44 $T=47840 29920 1 0 $X=47650 $Y=26960
X1591 VSS VDD 265 130 ICV_44 $T=47840 40800 1 0 $X=47650 $Y=37840
X1592 VSS VDD 228 178 ICV_44 $T=47840 100640 1 0 $X=47650 $Y=97680
X1593 VSS VDD 242 229 ICV_44 $T=47840 122400 1 0 $X=47650 $Y=119440
X1594 VSS VDD 341 396 ICV_44 $T=75900 127840 1 0 $X=75710 $Y=124880
X1595 VSS VDD 206 383 ICV_44 $T=75900 133280 1 0 $X=75710 $Y=130320
X1596 VSS VDD 413 392 ICV_44 $T=89700 40800 0 0 $X=89510 $Y=40560
X1597 VSS VDD 604 67 ICV_44 $T=117760 73440 0 0 $X=117570 $Y=73200
X1598 VSS VDD 604 140 ICV_44 $T=117760 89760 0 0 $X=117570 $Y=89520
X1599 VSS VDD 556 667 ICV_44 $T=117760 95200 0 0 $X=117570 $Y=94960
X1600 VSS VDD 343 602 ICV_44 $T=117760 122400 0 0 $X=117570 $Y=122160
X1601 VSS VDD 602 560 ICV_44 $T=117760 138720 0 0 $X=117570 $Y=138480
X1602 VSS VDD 67 563 ICV_44 $T=117760 144160 0 0 $X=117570 $Y=143920
X1603 VSS VDD 343 754 ICV_44 $T=132020 51680 1 0 $X=131830 $Y=48720
X1604 VSS VDD 510 387 ICV_44 $T=132020 73440 1 0 $X=131830 $Y=70480
X1605 VSS VDD 285 286 ICV_44 $T=132020 78880 1 0 $X=131830 $Y=75920
X1606 VSS VDD 109 116 152 135 ICV_45 $T=19780 84320 1 0 $X=19590 $Y=81360
X1607 VSS VDD 208 197 207 PAR_IN8<25> ICV_45 $T=33580 149600 0 0 $X=33390 $Y=149360
X1608 VSS VDD 442 420 293 PAR_IN3<21> ICV_45 $T=75900 24480 1 0 $X=75710 $Y=21520
X1609 VSS VDD 445 390 432 PAR_IN8<17> ICV_45 $T=75900 35360 1 0 $X=75710 $Y=32400
X1610 VSS VDD 449 486 513 PAR_IN7<7> ICV_45 $T=89700 149600 0 0 $X=89510 $Y=149360
X1611 VSS VDD 590 615 91 PAR_IN3<3> ICV_45 $T=103960 62560 1 0 $X=103770 $Y=59600
X1612 VSS VDD 659 693 289 PAR_IN3<19> ICV_45 $T=117760 78880 0 0 $X=117570 $Y=78640
X1613 VSS VDD 634 668 654 PAR_IN2<26> ICV_45 $T=117760 111520 0 0 $X=117570 $Y=111280
X1614 VSS VDD 121 644 677 PAR_IN7<12> ICV_45 $T=117760 133280 0 0 $X=117570 $Y=133040
X1615 VSS VDD 687 648 102 PAR_IN8<0> ICV_45 $T=117760 149600 0 0 $X=117570 $Y=149360
X1616 VSS VDD 731 765 654 PAR_IN2<18> ICV_45 $T=132020 68000 1 0 $X=131830 $Y=65040
X1617 VSS VDD ICV_46 $T=18400 155040 1 0 $X=18210 $Y=152080
X1618 VSS VDD ICV_46 $T=60260 73440 0 0 $X=60070 $Y=73200
X1619 VSS VDD ICV_46 $T=60260 127840 0 0 $X=60070 $Y=127600
X1620 VSS VDD ICV_46 $T=74520 29920 1 0 $X=74330 $Y=26960
X1621 VSS VDD ICV_46 $T=74520 62560 1 0 $X=74330 $Y=59600
X1622 VSS VDD ICV_46 $T=74520 73440 1 0 $X=74330 $Y=70480
X1623 VSS VDD ICV_46 $T=74520 138720 1 0 $X=74330 $Y=135760
X1624 VSS VDD ICV_46 $T=74520 144160 1 0 $X=74330 $Y=141200
X1625 VSS VDD ICV_46 $T=102580 35360 1 0 $X=102390 $Y=32400
X1626 VSS VDD ICV_46 $T=102580 84320 1 0 $X=102390 $Y=81360
X1627 VSS VDD ICV_46 $T=102580 116960 1 0 $X=102390 $Y=114000
X1628 VSS VDD ICV_46 $T=116380 68000 0 0 $X=116190 $Y=67760
X1629 VSS VDD ICV_46 $T=116380 100640 0 0 $X=116190 $Y=100400
X1630 VSS VDD ICV_46 $T=130640 19040 1 0 $X=130450 $Y=16080
X1631 VSS VDD ICV_46 $T=130640 111520 1 0 $X=130450 $Y=108560
X1632 VSS VDD ICV_46 $T=130640 116960 1 0 $X=130450 $Y=114000
X1633 VSS 119 ICV_47 $T=17940 89760 1 0 $X=17750 $Y=86800
X1634 VSS 116 ICV_47 $T=17940 95200 1 0 $X=17750 $Y=92240
X1635 VSS RESET ICV_47 $T=31740 19040 0 0 $X=31550 $Y=18800
X1636 VSS SERIAL_OUT ICV_47 $T=31740 24480 0 0 $X=31550 $Y=24240
X1637 VSS 201 ICV_47 $T=31740 62560 0 0 $X=31550 $Y=62320
X1638 VSS 203 ICV_47 $T=31740 122400 0 0 $X=31550 $Y=122160
X1639 VSS 180 ICV_47 $T=46000 73440 1 0 $X=45810 $Y=70480
X1640 VSS 37 ICV_47 $T=46000 78880 1 0 $X=45810 $Y=75920
X1641 VSS 316 ICV_47 $T=59800 19040 0 0 $X=59610 $Y=18800
X1642 VSS PAR_IN8<20> ICV_47 $T=59800 35360 0 0 $X=59610 $Y=35120
X1643 VSS 239 ICV_47 $T=59800 51680 0 0 $X=59610 $Y=51440
X1644 VSS 333 ICV_47 $T=59800 84320 0 0 $X=59610 $Y=84080
X1645 VSS 17 ICV_47 $T=59800 89760 0 0 $X=59610 $Y=89520
X1646 VSS PAR_IN7<14> ICV_47 $T=59800 106080 0 0 $X=59610 $Y=105840
X1647 VSS 336 ICV_47 $T=59800 133280 0 0 $X=59610 $Y=133040
X1648 VSS COUNT<4> ICV_47 $T=59800 138720 0 0 $X=59610 $Y=138480
X1649 VSS 420 ICV_47 $T=74060 19040 1 0 $X=73870 $Y=16080
X1650 VSS 423 ICV_47 $T=74060 95200 1 0 $X=73870 $Y=92240
X1651 VSS 352 ICV_47 $T=74060 100640 1 0 $X=73870 $Y=97680
X1652 VSS 336 ICV_47 $T=87860 19040 0 0 $X=87670 $Y=18800
X1653 VSS 81 ICV_47 $T=87860 95200 0 0 $X=87670 $Y=94960
X1654 VSS 500 ICV_47 $T=87860 106080 0 0 $X=87670 $Y=105840
X1655 VSS PAR_IN1<28> ICV_47 $T=87860 138720 0 0 $X=87670 $Y=138480
X1656 VSS 586 ICV_47 $T=102120 73440 1 0 $X=101930 $Y=70480
X1657 VSS PAR_IN5<27> ICV_47 $T=115920 29920 0 0 $X=115730 $Y=29680
X1658 VSS 510 ICV_47 $T=115920 40800 0 0 $X=115730 $Y=40560
X1659 VSS PAR_IN7<3> ICV_47 $T=115920 51680 0 0 $X=115730 $Y=51440
X1660 VSS PAR_IN6<1> ICV_47 $T=115920 127840 0 0 $X=115730 $Y=127600
X1661 VSS 695 ICV_47 $T=130180 29920 1 0 $X=129990 $Y=26960
X1662 VSS 728 ICV_47 $T=130180 57120 1 0 $X=129990 $Y=54160
X1663 VSS 628 ICV_47 $T=130180 122400 1 0 $X=129990 $Y=119440
X1664 VSS 736 ICV_47 $T=130180 127840 1 0 $X=129990 $Y=124880
X1665 VSS VDD ICV_48 $T=16100 19040 1 0 $X=15910 $Y=16080
X1666 VSS VDD ICV_48 $T=16100 73440 1 0 $X=15910 $Y=70480
X1667 VSS VDD ICV_48 $T=16100 149600 1 0 $X=15910 $Y=146640
X1668 VSS VDD ICV_48 $T=72220 84320 1 0 $X=72030 $Y=81360
X1669 VSS VDD ICV_48 $T=72220 111520 1 0 $X=72030 $Y=108560
X1670 VSS VDD ICV_48 $T=86020 29920 0 0 $X=85830 $Y=29680
X1671 VSS VDD ICV_48 $T=100280 29920 1 0 $X=100090 $Y=26960
X1672 VSS VDD ICV_48 $T=115920 13600 1 0 $X=115730 $Y=10640
X1673 VSS VDD ICV_48 $T=128340 40800 1 0 $X=128150 $Y=37840
X1674 VSS VDD 103 PAR_IN6<8> PAR_IN3<12> 128 158 178 PAR_IN3<12> ICV_49 $T=16560 133280 0 0 $X=16370 $Y=133040
X1675 VSS VDD 404 293 PAR_IN3<29> 426 421 293 PAR_IN3<29> ICV_49 $T=69460 35360 0 0 $X=69270 $Y=35120
X1676 VSS VDD 536 468 PAR_IN4<13> 256 468 431 PAR_IN4<13> ICV_49 $T=92920 84320 0 0 $X=92730 $Y=84080
X1677 VSS VDD 540 227 PAR_IN3<17> 579 581 91 PAR_IN3<17> ICV_49 $T=94300 57120 0 0 $X=94110 $Y=56880
X1678 VSS VDD 292 634 370 622 370 604 PAR_IN5<26> ICV_49 $T=109940 106080 1 0 $X=109750 $Y=103120
X1679 VSS VDD 343 625 PAR_IN6<6> 430 704 672 PAR_IN6<6> ICV_49 $T=121440 122400 0 0 $X=121250 $Y=122160
X1680 VSS VDD 696 510 PAR_IN3<2> 728 457 510 PAR_IN3<2> ICV_49 $T=121900 46240 0 0 $X=121710 $Y=46000
X1681 VSS VDD PAR_IN6<19> 513 PAR_IN7<23> 742 749 513 PAR_IN7<23> ICV_49 $T=125580 149600 0 0 $X=125390 $Y=149360
X1682 VSS VDD RESET 49 ICV_50 $T=7820 73440 1 0 $X=7630 $Y=70480
X1683 VSS VDD PAR_IN8<12> 87 ICV_50 $T=11040 127840 1 0 $X=10850 $Y=124880
X1684 VSS VDD PAR_IN5<7> 127 ICV_50 $T=20240 116960 0 0 $X=20050 $Y=116720
X1685 VSS VDD 145 176 ICV_50 $T=24380 13600 1 0 $X=24190 $Y=10640
X1686 VSS VDD 201 25 ICV_50 $T=37260 78880 0 0 $X=37070 $Y=78640
X1687 VSS VDD 228 231 ICV_50 $T=40020 13600 1 0 $X=39830 $Y=10640
X1688 VSS VDD 92 230 ICV_50 $T=40480 133280 0 0 $X=40290 $Y=133040
X1689 VSS VDD PAR_IN2<6> 290 ICV_50 $T=63020 84320 0 0 $X=62830 $Y=84080
X1690 VSS VDD 442 522 ICV_50 $T=92000 29920 1 0 $X=91810 $Y=26960
X1691 VSS VDD 169 494 ICV_50 $T=96140 24480 0 0 $X=95950 $Y=24240
X1692 VSS VDD 617 624 ICV_50 $T=107180 116960 1 0 $X=106990 $Y=114000
X1693 VSS VDD PAR_IN4<3> 181 ICV_50 $T=109480 46240 1 0 $X=109290 $Y=43280
X1694 VSS VDD 321 640 ICV_50 $T=109940 29920 1 0 $X=109750 $Y=26960
X1695 VSS VDD PAR_IN7<12> 644 ICV_50 $T=118680 133280 1 0 $X=118490 $Y=130320
X1696 VSS VDD 556 286 ICV_50 $T=121440 95200 0 0 $X=121250 $Y=94960
X1697 VSS VDD 301 677 ICV_50 $T=122820 106080 1 0 $X=122630 $Y=103120
X1698 VSS VDD PAR_IN5<7> 127 138 ICV_51 $T=19780 122400 1 0 $X=19590 $Y=119440
X1699 VSS VDD PAR_IN6<8> 103 129 ICV_51 $T=19780 138720 1 0 $X=19590 $Y=135760
X1700 VSS VDD COUNT<1> 34 246 ICV_51 $T=47840 95200 1 0 $X=47650 $Y=92240
X1701 VSS VDD PAR_IN2<12> 258 158 ICV_51 $T=47840 144160 1 0 $X=47650 $Y=141200
X1702 VSS VDD PAR_IN6<4> 103 244 ICV_51 $T=47840 155040 1 0 $X=47650 $Y=152080
X1703 VSS VDD PAR_IN6<28> 546 606 ICV_51 $T=103960 19040 1 0 $X=103770 $Y=16080
X1704 VSS VDD PAR_IN5<19> 563 619 ICV_51 $T=103960 46240 1 0 $X=103770 $Y=43280
X1705 VSS VDD PAR_IN2<8> 66 141 ICV_51 $T=103960 155040 1 0 $X=103770 $Y=152080
X1706 VSS VDD PAR_IN5<31> 127 629 ICV_51 $T=117760 13600 0 0 $X=117570 $Y=13360
X1707 VSS VDD PAR_IN5<1> 127 548 ICV_51 $T=117760 19040 0 0 $X=117570 $Y=18800
X1708 VSS VDD PAR_IN5<9> 620 389 ICV_51 $T=117760 24480 0 0 $X=117570 $Y=24240
X1709 VSS VDD PAR_IN6<13> 59 ICV_52 $T=7820 95200 1 0 $X=7630 $Y=92240
X1710 VSS VDD RESET 49 ICV_52 $T=7820 100640 1 0 $X=7630 $Y=97680
X1711 VSS VDD PAR_IN5<4> 67 ICV_52 $T=12880 13600 0 0 $X=12690 $Y=13360
X1712 VSS VDD PAR_IN2<5> 272 ICV_52 $T=49680 62560 0 0 $X=49490 $Y=62320
X1713 VSS VDD 375 393 ICV_52 $T=68080 62560 1 0 $X=67890 $Y=59600
X1714 VSS VDD 145 114 ICV_52 $T=78200 46240 1 0 $X=78010 $Y=43280
X1715 VSS VDD PAR_IN1<19> 401 ICV_52 $T=83260 13600 0 0 $X=83070 $Y=13360
X1716 VSS VDD 471 477 ICV_52 $T=84180 127840 1 0 $X=83990 $Y=124880
X1717 VSS VDD PAR_IN7<17> 127 ICV_52 $T=117300 19040 1 0 $X=117110 $Y=16080
X1718 VSS VDD 72 COUNT<0> ICV_53 $T=20240 46240 0 0 $X=20050 $Y=46000
X1719 VSS VDD 25 146 ICV_53 $T=20240 84320 0 0 $X=20050 $Y=84080
X1720 VSS VDD 282 334 ICV_53 $T=57500 78880 0 0 $X=57310 $Y=78640
X1721 VSS VDD 186 294 ICV_53 $T=58420 149600 1 0 $X=58230 $Y=146640
X1722 VSS VDD 373 392 ICV_53 $T=66240 51680 1 0 $X=66050 $Y=48720
X1723 VSS VDD 383 PAR_IN1<16> ICV_53 $T=76360 133280 0 0 $X=76170 $Y=133040
X1724 VSS VDD COUNT<4> 329 ICV_53 $T=78660 57120 0 0 $X=78470 $Y=56880
X1725 VSS VDD 280 468 ICV_53 $T=87400 24480 1 0 $X=87210 $Y=21520
X1726 VSS VDD 432 493 ICV_53 $T=99820 127840 1 0 $X=99630 $Y=124880
X1727 VSS VDD PAR_IN2<8> 67 ICV_53 $T=106720 149600 0 0 $X=106530 $Y=149360
X1728 VSS VDD PAR_IN5<23> 67 ICV_53 $T=113620 144160 0 0 $X=113430 $Y=143920
X1729 VSS VDD 113 COMPLETE VDD 116 VSS sky130_fd_sc_hd__or2_4 $T=15640 78880 0 0 $X=15450 $Y=78640
X1730 VSS VDD 186 PAR_IN1<12> VDD 195 VSS sky130_fd_sc_hd__or2_4 $T=28520 122400 1 0 $X=28330 $Y=119440
X1731 VSS VDD 193 146 VDD 152 VSS sky130_fd_sc_hd__or2_4 $T=30360 84320 1 0 $X=30170 $Y=81360
X1732 VSS VDD 206 PAR_IN1<10> VDD 217 VSS sky130_fd_sc_hd__or2_4 $T=34960 122400 0 0 $X=34770 $Y=122160
X1733 VSS VDD 206 PAR_IN1<26> VDD 219 VSS sky130_fd_sc_hd__or2_4 $T=34960 127840 0 0 $X=34770 $Y=127600
X1734 VSS VDD 186 PAR_IN1<8> VDD 224 VSS sky130_fd_sc_hd__or2_4 $T=35880 138720 1 0 $X=35690 $Y=135760
X1735 VSS VDD 25 201 VDD 13 VSS sky130_fd_sc_hd__or2_4 $T=37260 84320 1 0 $X=37070 $Y=81360
X1736 VSS VDD 222 229 VDD 193 VSS sky130_fd_sc_hd__or2_4 $T=39560 84320 0 0 $X=39370 $Y=84080
X1737 VSS VDD 13 18 VDD 222 VSS sky130_fd_sc_hd__or2_4 $T=40940 95200 0 0 $X=40750 $Y=94960
X1738 VSS VDD 281 PAR_IN1<24> VDD 308 VSS sky130_fd_sc_hd__or2_4 $T=53360 122400 1 0 $X=53170 $Y=119440
X1739 VSS VDD 281 PAR_IN1<9> VDD 309 VSS sky130_fd_sc_hd__or2_4 $T=53360 127840 0 0 $X=53170 $Y=127600
X1740 VSS VDD 303 PAR_IN1<18> VDD 317 VSS sky130_fd_sc_hd__or2_4 $T=54740 62560 1 0 $X=54550 $Y=59600
X1741 VSS VDD 303 PAR_IN1<2> VDD 326 VSS sky130_fd_sc_hd__or2_4 $T=56580 68000 1 0 $X=56390 $Y=65040
X1742 VSS VDD 186 PAR_IN1<4> VDD 283 VSS sky130_fd_sc_hd__or2_4 $T=57500 155040 1 0 $X=57310 $Y=152080
X1743 VSS VDD 300 SAMPLE_COUNT<3> VDD 340 VSS sky130_fd_sc_hd__or2_4 $T=58880 51680 1 0 $X=58690 $Y=48720
X1744 VSS VDD 303 PAR_IN1<14> VDD 393 VSS sky130_fd_sc_hd__or2_4 $T=66240 57120 1 0 $X=66050 $Y=54160
X1745 VSS VDD 392 PAR_IN1<13> VDD 394 VSS sky130_fd_sc_hd__or2_4 $T=68540 51680 0 0 $X=68350 $Y=51440
X1746 VSS VDD 401 PAR_IN1<7> VDD 410 VSS sky130_fd_sc_hd__or2_4 $T=69000 84320 1 0 $X=68810 $Y=81360
X1747 VSS VDD 385 COUNT<1> VDD 21 VSS sky130_fd_sc_hd__or2_4 $T=69460 95200 0 0 $X=69270 $Y=94960
X1748 VSS VDD 413 PAR_IN1<20> VDD 418 VSS sky130_fd_sc_hd__or2_4 $T=75900 13600 0 0 $X=75710 $Y=13360
X1749 VSS VDD 401 PAR_IN1<31> VDD 455 VSS sky130_fd_sc_hd__or2_4 $T=77280 19040 1 0 $X=77090 $Y=16080
X1750 VSS VDD 401 PAR_IN1<23> VDD 456 VSS sky130_fd_sc_hd__or2_4 $T=77280 111520 1 0 $X=77090 $Y=108560
X1751 VSS VDD 186 PAR_IN1<25> VDD 406 VSS sky130_fd_sc_hd__or2_4 $T=79580 144160 0 0 $X=79390 $Y=143920
X1752 VSS VDD 413 PAR_IN1<15> VDD 478 VSS sky130_fd_sc_hd__or2_4 $T=80500 133280 0 0 $X=80310 $Y=133040
X1753 VSS VDD 281 PAR_IN1<16> VDD 467 VSS sky130_fd_sc_hd__or2_4 $T=81880 138720 1 0 $X=81690 $Y=135760
X1754 VSS VDD 392 PAR_IN1<11> VDD 487 VSS sky130_fd_sc_hd__or2_4 $T=82340 78880 0 0 $X=82150 $Y=78640
X1755 VSS VDD 401 PAR_IN1<19> VDD 489 VSS sky130_fd_sc_hd__or2_4 $T=83260 19040 1 0 $X=83070 $Y=16080
X1756 VSS VDD 383 PAR_IN1<0> VDD 451 VSS sky130_fd_sc_hd__or2_4 $T=83260 149600 1 0 $X=83070 $Y=146640
X1757 VSS VDD 303 PAR_IN1<22> VDD 481 VSS sky130_fd_sc_hd__or2_4 $T=83720 122400 1 0 $X=83530 $Y=119440
X1758 VSS VDD 303 PAR_IN1<30> VDD 433 VSS sky130_fd_sc_hd__or2_4 $T=87860 57120 1 0 $X=87670 $Y=54160
X1759 VSS VDD 186 PAR_IN1<1> VDD 500 VSS sky130_fd_sc_hd__or2_4 $T=91080 111520 0 0 $X=90890 $Y=111280
X1760 VSS VDD 281 PAR_IN1<28> VDD 472 VSS sky130_fd_sc_hd__or2_4 $T=91080 138720 0 0 $X=90890 $Y=138480
X1761 VSS VDD 413 PAR_IN1<17> VDD 526 VSS sky130_fd_sc_hd__or2_4 $T=92000 13600 0 0 $X=91810 $Y=13360
X1762 VSS VDD 401 PAR_IN1<27> VDD 543 VSS sky130_fd_sc_hd__or2_4 $T=94300 19040 1 0 $X=94110 $Y=16080
X1763 VSS VDD 392 PAR_IN1<29> VDD 490 VSS sky130_fd_sc_hd__or2_4 $T=99360 29920 0 0 $X=99170 $Y=29680
X1764 VSS VDD 413 PAR_IN1<3> VDD 540 VSS sky130_fd_sc_hd__or2_4 $T=99820 13600 0 0 $X=99630 $Y=13360
X1765 VSS VDD 392 PAR_IN1<5> VDD 535 VSS sky130_fd_sc_hd__or2_4 $T=100740 78880 0 0 $X=100550 $Y=78640
X1766 VSS VDD 392 PAR_IN1<21> VDD 523 VSS sky130_fd_sc_hd__or2_4 $T=106260 29920 0 0 $X=106070 $Y=29680
X1767 VSS VDD ICV_54 $T=19780 100640 1 0 $X=19590 $Y=97680
X1768 VSS VDD ICV_54 $T=47840 68000 1 0 $X=47650 $Y=65040
X1769 VSS VDD ICV_54 $T=47840 138720 1 0 $X=47650 $Y=135760
X1770 VSS VDD ICV_54 $T=61640 116960 0 0 $X=61450 $Y=116720
X1771 VSS VDD ICV_54 $T=61640 144160 0 0 $X=61450 $Y=143920
X1772 VSS VDD ICV_54 $T=89700 35360 0 0 $X=89510 $Y=35120
X1773 VSS VDD ICV_54 $T=103960 68000 1 0 $X=103770 $Y=65040
X1774 VSS VDD ICV_54 $T=103960 144160 1 0 $X=103770 $Y=141200
X1775 VSS VDD 203 195 163 VDD 218 VSS sky130_fd_sc_hd__and3_4 $T=34040 127840 1 0 $X=33850 $Y=124880
X1776 VSS VDD 227 224 196 VDD 243 VSS sky130_fd_sc_hd__and3_4 $T=40020 133280 1 0 $X=39830 $Y=130320
X1777 VSS VDD 262 217 274 VDD 259 VSS sky130_fd_sc_hd__and3_4 $T=48760 116960 0 0 $X=48570 $Y=116720
X1778 VSS VDD 203 309 323 VDD 358 VSS sky130_fd_sc_hd__and3_4 $T=60720 133280 1 0 $X=60530 $Y=130320
X1779 VSS VDD 262 326 320 VDD 337 VSS sky130_fd_sc_hd__and3_4 $T=61180 73440 1 0 $X=60990 $Y=70480
X1780 VSS VDD 135 394 287 VDD 409 VSS sky130_fd_sc_hd__and3_4 $T=68080 73440 0 0 $X=67890 $Y=73200
X1781 VSS VDD 396 406 214 VDD 397 VSS sky130_fd_sc_hd__and3_4 $T=69920 138720 0 0 $X=69730 $Y=138480
X1782 VSS VDD COUNT<4> 433 416 VDD 375 VSS sky130_fd_sc_hd__and3_4 $T=77280 62560 1 0 $X=77090 $Y=59600
X1783 VSS VDD 203 451 453 VDD 412 VSS sky130_fd_sc_hd__and3_4 $T=77740 144160 1 0 $X=77550 $Y=141200
X1784 VSS VDD 396 455 474 VDD 482 VSS sky130_fd_sc_hd__and3_4 $T=81880 29920 0 0 $X=81690 $Y=29680
X1785 VSS VDD 341 472 477 VDD 253 VSS sky130_fd_sc_hd__and3_4 $T=81880 127840 0 0 $X=81690 $Y=127600
X1786 VSS VDD 341 481 450 VDD 379 VSS sky130_fd_sc_hd__and3_4 $T=82800 116960 1 0 $X=82610 $Y=114000
X1787 VSS VDD 469 490 458 VDD 408 VSS sky130_fd_sc_hd__and3_4 $T=85100 40800 1 0 $X=84910 $Y=37840
X1788 VSS VDD 227 500 512 VDD 476 VSS sky130_fd_sc_hd__and3_4 $T=89240 111520 1 0 $X=89050 $Y=108560
X1789 VSS VDD 135 487 517 VDD 497 VSS sky130_fd_sc_hd__and3_4 $T=90160 78880 1 0 $X=89970 $Y=75920
X1790 VSS VDD 469 523 525 VDD 495 VSS sky130_fd_sc_hd__and3_4 $T=91080 35360 1 0 $X=90890 $Y=32400
X1791 VSS VDD 227 478 530 VDD 483 VSS sky130_fd_sc_hd__and3_4 $T=91080 127840 0 0 $X=90890 $Y=127600
X1792 VSS VDD 396 526 509 VDD 506 VSS sky130_fd_sc_hd__and3_4 $T=91540 35360 0 0 $X=91350 $Y=35120
X1793 VSS VDD 135 535 536 VDD 505 VSS sky130_fd_sc_hd__and3_4 $T=92920 78880 0 0 $X=92730 $Y=78640
X1794 VSS VDD 469 543 549 VDD 527 VSS sky130_fd_sc_hd__and3_4 $T=95680 40800 1 0 $X=95490 $Y=37840
X1795 VSS VDD 210 211 184 12 115 ICV_55 $T=34960 46240 0 0 $X=34770 $Y=46000
X1796 VSS VDD COUNT<4> COUNT<4> 219 237 248 ICV_55 $T=40940 116960 0 0 $X=40750 $Y=116720
X1797 VSS VDD 268 240 265 268 300 ICV_55 $T=51060 46240 1 0 $X=50870 $Y=43280
X1798 VSS VDD 245 203 283 245 305 ICV_55 $T=51520 138720 0 0 $X=51330 $Y=138480
X1799 VSS VDD 358 341 308 335 257 ICV_55 $T=61640 127840 1 0 $X=61450 $Y=124880
X1800 VSS VDD 357 COUNT<4> 317 357 334 ICV_55 $T=63020 68000 0 0 $X=62830 $Y=67760
X1801 VSS VDD 400 262 393 400 356 ICV_55 $T=67620 62560 0 0 $X=67430 $Y=62320
X1802 VSS VDD PAR_IN8<17> 396 418 377 306 ICV_55 $T=73600 29920 0 0 $X=73410 $Y=29680
X1803 VSS VDD 460 227 410 447 460 ICV_55 $T=77280 95200 1 0 $X=77090 $Y=92240
X1804 VSS VDD 467 341 467 471 382 ICV_55 $T=81420 122400 0 0 $X=81230 $Y=122160
X1805 VSS VDD 506 469 456 492 448 ICV_55 $T=85100 95200 1 0 $X=84910 $Y=92240
X1806 VSS VDD 534 469 489 534 491 ICV_55 $T=92000 62560 0 0 $X=91810 $Y=62320
X1807 VSS VDD 581 227 540 550 511 ICV_55 $T=96140 62560 1 0 $X=95950 $Y=59600
X1808 VSS VDD 191 82 157 VDD 204 VSS sky130_fd_sc_hd__nor3_4 $T=27600 46240 1 0 $X=27410 $Y=43280
X1809 VSS VDD COUNT<0> 246 247 VDD 223 VSS sky130_fd_sc_hd__nor3_4 $T=44160 89760 0 0 $X=43970 $Y=89520
X1810 VSS VDD 229 253 218 VDD 252 VSS sky130_fd_sc_hd__nor3_4 $T=49220 127840 1 0 $X=49030 $Y=124880
X1811 VSS VDD 14 252 278 VDD 291 VSS sky130_fd_sc_hd__nor3_4 $T=49680 106080 0 0 $X=49490 $Y=105840
X1812 VSS VDD 118 257 243 VDD 313 VSS sky130_fd_sc_hd__nor3_4 $T=51520 122400 0 0 $X=51330 $Y=122160
X1813 VSS VDD COUNT<2> 312 313 VDD 279 VSS sky130_fd_sc_hd__nor3_4 $T=54740 116960 1 0 $X=54550 $Y=114000
X1814 VSS VDD 319 305 306 VDD 278 VSS sky130_fd_sc_hd__nor3_4 $T=57040 111520 1 0 $X=56850 $Y=108560
X1815 VSS VDD 229 358 397 VDD 403 VSS sky130_fd_sc_hd__nor3_4 $T=64400 127840 0 0 $X=64210 $Y=127600
X1816 VSS VDD COUNT<2> 403 365 VDD 385 VSS sky130_fd_sc_hd__nor3_4 $T=69000 100640 0 0 $X=68810 $Y=100400
X1817 VSS VDD 319 412 382 VDD 312 VSS sky130_fd_sc_hd__nor3_4 $T=70840 122400 0 0 $X=70650 $Y=122160
X1818 VSS VDD 118 408 409 VDD 434 VSS sky130_fd_sc_hd__nor3_4 $T=74980 68000 0 0 $X=74790 $Y=67760
X1819 VSS VDD 14 411 436 VDD 24 VSS sky130_fd_sc_hd__nor3_4 $T=74980 84320 0 0 $X=74790 $Y=84080
X1820 VSS VDD 14 422 434 VDD 22 VSS sky130_fd_sc_hd__nor3_4 $T=77280 78880 1 0 $X=77090 $Y=75920
X1821 VSS VDD 202 460 448 VDD 436 VSS sky130_fd_sc_hd__nor3_4 $T=78200 89760 0 0 $X=78010 $Y=89520
X1822 VSS VDD 118 483 482 VDD 411 VSS sky130_fd_sc_hd__nor3_4 $T=81420 89760 1 0 $X=81230 $Y=86800
X1823 VSS VDD COUNT<2> 488 479 VDD 23 VSS sky130_fd_sc_hd__nor3_4 $T=83260 73440 1 0 $X=83070 $Y=70480
X1824 VSS VDD 202 476 506 VDD 365 VSS sky130_fd_sc_hd__nor3_4 $T=84640 100640 1 0 $X=84450 $Y=97680
X1825 VSS VDD 202 511 491 VDD 488 VSS sky130_fd_sc_hd__nor3_4 $T=89240 68000 1 0 $X=89050 $Y=65040
X1826 VSS VDD 118 527 497 VDD 479 VSS sky130_fd_sc_hd__nor3_4 $T=91080 68000 0 0 $X=90890 $Y=67760
X1827 VSS VDD 202 505 495 VDD 422 VSS sky130_fd_sc_hd__nor3_4 $T=91080 73440 0 0 $X=90890 $Y=73200
X1828 VSS VDD COMPLETE VDD 72 VSS sky130_fd_sc_hd__inv_8 $T=10120 51680 1 0 $X=9930 $Y=48720
X1829 VSS VDD INTERNAL_FINISH VDD 5 VSS sky130_fd_sc_hd__inv_8 $T=10120 68000 0 0 $X=9930 $Y=67760
X1830 VSS VDD 83 VDD 113 VSS sky130_fd_sc_hd__inv_8 $T=14260 62560 0 0 $X=14070 $Y=62320
X1831 VSS VDD COUNT<1> VDD 25 VSS sky130_fd_sc_hd__inv_8 $T=25300 106080 1 0 $X=25110 $Y=103120
X1832 VSS VDD 133 VDD 12 VSS sky130_fd_sc_hd__inv_8 $T=25760 68000 0 0 $X=25570 $Y=67760
X1833 VSS VDD COUNT<5> VDD 194 VSS sky130_fd_sc_hd__inv_8 $T=27140 73440 1 0 $X=26950 $Y=70480
X1834 VSS VDD COUNT<0> VDD 201 VSS sky130_fd_sc_hd__inv_8 $T=34960 73440 1 0 $X=34770 $Y=70480
X1835 VSS VDD 222 VDD 11 VSS sky130_fd_sc_hd__inv_8 $T=37720 95200 1 0 $X=37530 $Y=92240
X1836 VSS VDD SAMPLE_COUNT<3> VDD 239 VSS sky130_fd_sc_hd__inv_8 $T=40020 46240 1 0 $X=39830 $Y=43280
X1837 VSS VDD COUNT<3> VDD 242 VSS sky130_fd_sc_hd__inv_8 $T=40020 122400 1 0 $X=39830 $Y=119440
X1838 VSS VDD SAMPLE_COUNT<2> VDD 268 VSS sky130_fd_sc_hd__inv_8 $T=46460 51680 0 0 $X=46270 $Y=51440
X1839 VSS VDD COUNT<2> VDD 18 VSS sky130_fd_sc_hd__inv_8 $T=48760 95200 0 0 $X=48570 $Y=94960
X1840 VSS VDD SAMPLE_COUNT<1> VDD 240 VSS sky130_fd_sc_hd__inv_8 $T=49220 35360 1 0 $X=49030 $Y=32400
X1841 VSS VDD SAMPLE_COUNT<0> VDD 265 VSS sky130_fd_sc_hd__inv_8 $T=49680 35360 0 0 $X=49490 $Y=35120
X1842 VSS VDD COUNT<4> VDD 351 VSS sky130_fd_sc_hd__inv_8 $T=60260 144160 1 0 $X=60070 $Y=141200
X1843 VSS VDD 457 VDD 206 VSS sky130_fd_sc_hd__inv_8 $T=81880 111520 0 0 $X=81690 $Y=111280
X1844 VSS VDD 83 97 76 VDD 75 VSS sky130_fd_sc_hd__o21a_4 $T=10580 35360 1 0 $X=10390 $Y=32400
X1845 VSS VDD READY 69 5 VDD 83 VSS sky130_fd_sc_hd__o21a_4 $T=10580 62560 1 0 $X=10390 $Y=59600
X1846 VSS VDD 130 6 7 VDD 157 VSS sky130_fd_sc_hd__o21a_4 $T=24380 46240 0 0 $X=24190 $Y=46000
X1847 VSS VDD 13 COUNT<0> COUNT<1> VDD 119 VSS sky130_fd_sc_hd__o21a_4 $T=28520 95200 1 0 $X=28330 $Y=92240
X1848 VSS VDD 201 146 COUNT<5> VDD 192 VSS sky130_fd_sc_hd__o21a_4 $T=31280 68000 1 0 $X=31090 $Y=65040
X1849 VSS VDD 193 202 11 VDD 136 VSS sky130_fd_sc_hd__o21a_4 $T=34500 89760 1 0 $X=34310 $Y=86800
X1850 VSS VDD 143 130 133 VDD 210 VSS sky130_fd_sc_hd__o21a_4 $T=34960 51680 0 0 $X=34770 $Y=51440
X1851 VSS VDD 194 135 193 VDD 166 VSS sky130_fd_sc_hd__o21a_4 $T=34960 78880 1 0 $X=34770 $Y=75920
X1852 VSS VDD 25 279 291 VDD 247 VSS sky130_fd_sc_hd__o21a_4 $T=49220 106080 1 0 $X=49030 $Y=103120
X1853 VSS VDD 351 PAR_IN1<6> 383 VDD 353 VSS sky130_fd_sc_hd__o21a_4 $T=63480 144160 0 0 $X=63290 $Y=143920
X1854 VSS VDD COUNT<2> 379 361 VDD 20 VSS sky130_fd_sc_hd__o21a_4 $T=66700 111520 1 0 $X=66510 $Y=108560
X1855 VSS VDD 210 115 146 VDD 198 VSS sky130_fd_sc_hd__or3_4 $T=35880 57120 1 0 $X=35690 $Y=54160
X1856 VSS VDD 248 259 242 VDD 17 VSS sky130_fd_sc_hd__or3_4 $T=47380 111520 0 0 $X=47190 $Y=111280
X1857 VSS VDD 337 334 319 VDD 16 VSS sky130_fd_sc_hd__or3_4 $T=60720 84320 1 0 $X=60530 $Y=81360
X1858 VSS VDD 356 375 229 VDD 19 VSS sky130_fd_sc_hd__or3_4 $T=66240 68000 1 0 $X=66050 $Y=65040
X1859 VSS VDD 97 4 COUNT<5> 83 VDD 105 VSS sky130_fd_sc_hd__and4_4 $T=21160 29920 1 0 $X=20970 $Y=26960
X1860 VSS VDD 100 56 READY 64 VDD 98 VSS sky130_fd_sc_hd__and4_4 $T=21160 62560 1 0 $X=20970 $Y=59600
X1861 VSS VDD 184 12 69 4 VDD 191 VSS sky130_fd_sc_hd__and4_4 $T=28060 57120 1 0 $X=27870 $Y=54160
X1862 VSS VDD 215 56 143 130 VDD 271 VSS sky130_fd_sc_hd__and4_4 $T=46460 46240 0 0 $X=46270 $Y=46000
X1863 VSS VDD 239 SAMPLE_COUNT<2> 143 184 VDD 264 VSS sky130_fd_sc_hd__and4_4 $T=46920 40800 0 0 $X=46730 $Y=40560
X1864 VSS VDD 215 268 143 184 VDD 282 VSS sky130_fd_sc_hd__and4_4 $T=48760 57120 0 0 $X=48570 $Y=56880
X1865 VSS VDD 215 56 211 130 VDD 285 VSS sky130_fd_sc_hd__and4_4 $T=49220 57120 1 0 $X=49030 $Y=54160
X1866 VSS VDD 215 268 211 130 VDD 301 VSS sky130_fd_sc_hd__and4_4 $T=51060 51680 1 0 $X=50870 $Y=48720
X1867 VSS VDD 211 184 239 SAMPLE_COUNT<2> VDD 329 VSS sky130_fd_sc_hd__and4_4 $T=56120 57120 1 0 $X=55930 $Y=54160
X1868 VSS VDD 211 SAMPLE_COUNT<0> 239 268 VDD 343 VSS sky130_fd_sc_hd__and4_4 $T=58880 46240 1 0 $X=58690 $Y=43280
X1869 VSS VDD 56 64 VDD 65 VSS sky130_fd_sc_hd__nor2_4 $T=10120 40800 1 0 $X=9930 $Y=37840
X1870 VSS VDD 82 26 VDD 58 VSS sky130_fd_sc_hd__nor2_4 $T=10120 57120 1 0 $X=9930 $Y=54160
X1871 VSS VDD 232 234 VDD 205 VSS sky130_fd_sc_hd__nor2_4 $T=40480 68000 0 0 $X=40290 $Y=67760
X1872 VSS VDD 49 55 RESET VDD SAMPLE_COUNT<2> VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 29920 0 0 $X=7630 $Y=29680
X1873 VSS VDD 49 58 RESET VDD INTERNAL_FINISH VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 73440 0 0 $X=7630 $Y=73200
X1874 VSS VDD 49 60 RESET VDD COUNT<4> VSS sky130_fd_sc_hd__dfrtp_4 $T=7820 100640 0 0 $X=7630 $Y=100400
X1875 VSS VDD 49 98 RESET VDD COMPLETE VSS sky130_fd_sc_hd__dfrtp_4 $T=11500 57120 0 0 $X=11310 $Y=56880
X1876 VSS VDD 49 105 RESET VDD COUNT<5> VSS sky130_fd_sc_hd__dfrtp_4 $T=13340 19040 0 0 $X=13150 $Y=18800
X1877 VSS VDD 49 75 RESET VDD SAMPLE_COUNT<3> VSS sky130_fd_sc_hd__dfrtp_4 $T=13340 35360 0 0 $X=13150 $Y=35120
X1878 VSS VDD 49 110 RESET VDD COUNT<1> VSS sky130_fd_sc_hd__dfrtp_4 $T=14720 106080 0 0 $X=14530 $Y=105840
X1879 VSS VDD 165 177 RESET VDD SERIAL_OUT VSS sky130_fd_sc_hd__dfrtp_4 $T=25300 24480 1 0 $X=25110 $Y=21520
X1880 VSS VDD 165 174 RESET VDD COUNT<0> VSS sky130_fd_sc_hd__dfrtp_4 $T=25760 35360 1 0 $X=25570 $Y=32400
X1881 VSS VDD 165 167 RESET VDD COUNT<3> VSS sky130_fd_sc_hd__dfrtp_4 $T=27600 111520 1 0 $X=27410 $Y=108560
X1882 VSS VDD 165 171 RESET VDD COUNT<2> VSS sky130_fd_sc_hd__dfrtp_4 $T=33120 106080 1 0 $X=32930 $Y=103120
X1883 VSS VDD 165 190 RESET VDD SAMPLE_COUNT<1> VSS sky130_fd_sc_hd__dfrtp_4 $T=34960 19040 0 0 $X=34770 $Y=18800
X1884 VSS VDD 165 204 RESET VDD SAMPLE_COUNT<0> VSS sky130_fd_sc_hd__dfrtp_4 $T=34960 29920 0 0 $X=34770 $Y=29680
X1885 VSS VDD 29 49 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=11040 62560 0 0 $X=10850 $Y=62320
X1886 VSS VDD 29 165 VDD VSS sky130_fd_sc_hd__clkbuf_1 $T=28980 57120 0 0 $X=28790 $Y=56880
X1887 VSS VDD 109 12 100 60 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=14260 89760 0 0 $X=14070 $Y=89520
X1888 VSS VDD 108 107 100 110 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=14260 95200 0 0 $X=14070 $Y=94960
X1889 VSS VDD 155 183 100 167 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=23920 100640 0 0 $X=23730 $Y=100400
X1890 VSS VDD 154 30 100 171 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=25300 100640 1 0 $X=25110 $Y=97680
X1891 VSS VDD 170 198 4 190 VDD VSS sky130_fd_sc_hd__a21oi_4 $T=27600 40800 1 0 $X=27410 $Y=37840
X1892 VSS VDD 119 133 VDD 107 VSS sky130_fd_sc_hd__nand2_4 $T=21160 95200 1 0 $X=20970 $Y=92240
X1893 VSS VDD 136 133 VDD 183 VSS sky130_fd_sc_hd__nand2_4 $T=25760 95200 0 0 $X=25570 $Y=94960
X1894 VSS VDD 76 65 82 97 4 55 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=8740 40800 0 0 $X=8550 $Y=40560
X1895 VSS VDD 82 6 192 69 COUNT<0> 174 VDD VSS sky130_fd_sc_hd__a2111oi_4 $T=24840 51680 1 0 $X=24650 $Y=48720
X1896 VSS VDD ICV_56 $T=5520 51680 0 0 $X=5330 $Y=51440
X1897 VSS VDD ICV_56 $T=5520 106080 0 0 $X=5330 $Y=105840
X1898 VSS VDD ICV_56 $T=5520 111520 1 0 $X=5330 $Y=108560
X1899 VSS VDD ICV_56 $T=5520 122400 1 0 $X=5330 $Y=119440
X1900 VSS VDD ICV_56 $T=5520 122400 0 0 $X=5330 $Y=122160
X1901 VSS VDD ICV_56 $T=5520 127840 1 0 $X=5330 $Y=124880
X1902 VSS VDD ICV_56 $T=5520 127840 0 0 $X=5330 $Y=127600
X1903 VSS VDD ICV_56 $T=5520 133280 1 0 $X=5330 $Y=130320
.ENDS
***************************************
