VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

MACRO deserialiser_unit_cell_1
  CLASS BLOCK ;
  FOREIGN deserialiser_unit_cell_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 356.165 BY 366.885 ;
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END CLK
  PIN COMPLETE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 362.885 66.150 366.885 ;
    END
  END COMPLETE
  PIN COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END COUNT[0]
  PIN COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 254.360 356.165 254.960 ;
    END
  END COUNT[1]
  PIN COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 25.200 356.165 25.800 ;
    END
  END COUNT[2]
  PIN COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 362.885 248.770 366.885 ;
    END
  END COUNT[3]
  PIN COUNT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.830 362.885 78.110 366.885 ;
    END
  END COUNT[4]
  PIN COUNT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END COUNT[5]
  PIN INTERNAL_FINISH
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.050 362.885 58.330 366.885 ;
    END
  END INTERNAL_FINISH
  PIN OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.070 362.885 328.350 366.885 ;
    END
  END OUT[0]
  PIN OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 362.885 125.490 366.885 ;
    END
  END OUT[10]
  PIN OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.450 362.885 145.730 366.885 ;
    END
  END OUT[11]
  PIN OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END OUT[12]
  PIN OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END OUT[13]
  PIN OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END OUT[14]
  PIN OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 362.885 133.770 366.885 ;
    END
  END OUT[15]
  PIN OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 272.410 362.885 272.690 366.885 ;
    END
  END OUT[16]
  PIN OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END OUT[17]
  PIN OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END OUT[18]
  PIN OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END OUT[19]
  PIN OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END OUT[1]
  PIN OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END OUT[20]
  PIN OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END OUT[21]
  PIN OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.030 362.885 340.310 366.885 ;
    END
  END OUT[22]
  PIN OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 362.885 105.710 366.885 ;
    END
  END OUT[23]
  PIN OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END OUT[24]
  PIN OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 284.370 362.885 284.650 366.885 ;
    END
  END OUT[25]
  PIN OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 362.885 81.790 366.885 ;
    END
  END OUT[26]
  PIN OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END OUT[27]
  PIN OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END OUT[28]
  PIN OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END OUT[29]
  PIN OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END OUT[2]
  PIN OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END OUT[30]
  PIN OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END OUT[31]
  PIN OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END OUT[3]
  PIN OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END OUT[4]
  PIN OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 213.560 356.165 214.160 ;
    END
  END OUT[5]
  PIN OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 362.885 97.890 366.885 ;
    END
  END OUT[6]
  PIN OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END OUT[7]
  PIN OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END OUT[8]
  PIN OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 362.885 34.410 366.885 ;
    END
  END OUT[9]
  PIN PAR_IN1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 331.200 356.165 331.800 ;
    END
  END PAR_IN1[0]
  PIN PAR_IN1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 160.520 356.165 161.120 ;
    END
  END PAR_IN1[10]
  PIN PAR_IN1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END PAR_IN1[11]
  PIN PAR_IN1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.070 362.885 213.350 366.885 ;
    END
  END PAR_IN1[12]
  PIN PAR_IN1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END PAR_IN1[13]
  PIN PAR_IN1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 362.885 42.230 366.885 ;
    END
  END PAR_IN1[14]
  PIN PAR_IN1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 231.240 356.165 231.840 ;
    END
  END PAR_IN1[15]
  PIN PAR_IN1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END PAR_IN1[16]
  PIN PAR_IN1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END PAR_IN1[17]
  PIN PAR_IN1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END PAR_IN1[18]
  PIN PAR_IN1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 131.280 356.165 131.880 ;
    END
  END PAR_IN1[19]
  PIN PAR_IN1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 362.885 46.370 366.885 ;
    END
  END PAR_IN1[1]
  PIN PAR_IN1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END PAR_IN1[20]
  PIN PAR_IN1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END PAR_IN1[21]
  PIN PAR_IN1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 260.480 356.165 261.080 ;
    END
  END PAR_IN1[22]
  PIN PAR_IN1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 102.040 356.165 102.640 ;
    END
  END PAR_IN1[23]
  PIN PAR_IN1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.790 362.885 205.070 366.885 ;
    END
  END PAR_IN1[24]
  PIN PAR_IN1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.750 362.885 102.030 366.885 ;
    END
  END PAR_IN1[25]
  PIN PAR_IN1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.250 362.885 320.530 366.885 ;
    END
  END PAR_IN1[26]
  PIN PAR_IN1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 207.440 356.165 208.040 ;
    END
  END PAR_IN1[27]
  PIN PAR_IN1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END PAR_IN1[28]
  PIN PAR_IN1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 42.880 356.165 43.480 ;
    END
  END PAR_IN1[29]
  PIN PAR_IN1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 125.160 356.165 125.760 ;
    END
  END PAR_IN1[2]
  PIN PAR_IN1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 362.885 121.810 366.885 ;
    END
  END PAR_IN1[30]
  PIN PAR_IN1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END PAR_IN1[31]
  PIN PAR_IN1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 31.320 356.165 31.920 ;
    END
  END PAR_IN1[3]
  PIN PAR_IN1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END PAR_IN1[4]
  PIN PAR_IN1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END PAR_IN1[5]
  PIN PAR_IN1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END PAR_IN1[6]
  PIN PAR_IN1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END PAR_IN1[7]
  PIN PAR_IN1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.850 362.885 348.130 366.885 ;
    END
  END PAR_IN1[8]
  PIN PAR_IN1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END PAR_IN1[9]
  PIN PAR_IN2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END PAR_IN2[0]
  PIN PAR_IN2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 362.885 6.350 366.885 ;
    END
  END PAR_IN2[10]
  PIN PAR_IN2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END PAR_IN2[11]
  PIN PAR_IN2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END PAR_IN2[12]
  PIN PAR_IN2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END PAR_IN2[13]
  PIN PAR_IN2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END PAR_IN2[14]
  PIN PAR_IN2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 202.000 356.165 202.600 ;
    END
  END PAR_IN2[15]
  PIN PAR_IN2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 236.680 356.165 237.280 ;
    END
  END PAR_IN2[16]
  PIN PAR_IN2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END PAR_IN2[17]
  PIN PAR_IN2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END PAR_IN2[18]
  PIN PAR_IN2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 256.770 362.885 257.050 366.885 ;
    END
  END PAR_IN2[19]
  PIN PAR_IN2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END PAR_IN2[1]
  PIN PAR_IN2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END PAR_IN2[20]
  PIN PAR_IN2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END PAR_IN2[21]
  PIN PAR_IN2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.350 362.885 14.630 366.885 ;
    END
  END PAR_IN2[22]
  PIN PAR_IN2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 60.560 356.165 61.160 ;
    END
  END PAR_IN2[23]
  PIN PAR_IN2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END PAR_IN2[24]
  PIN PAR_IN2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END PAR_IN2[25]
  PIN PAR_IN2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 325.080 356.165 325.680 ;
    END
  END PAR_IN2[26]
  PIN PAR_IN2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END PAR_IN2[27]
  PIN PAR_IN2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 242.800 356.165 243.400 ;
    END
  END PAR_IN2[28]
  PIN PAR_IN2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END PAR_IN2[29]
  PIN PAR_IN2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END PAR_IN2[2]
  PIN PAR_IN2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END PAR_IN2[30]
  PIN PAR_IN2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END PAR_IN2[31]
  PIN PAR_IN2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END PAR_IN2[3]
  PIN PAR_IN2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.830 362.885 193.110 366.885 ;
    END
  END PAR_IN2[4]
  PIN PAR_IN2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.050 362.885 173.330 366.885 ;
    END
  END PAR_IN2[5]
  PIN PAR_IN2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END PAR_IN2[6]
  PIN PAR_IN2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END PAR_IN2[7]
  PIN PAR_IN2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 362.885 129.630 366.885 ;
    END
  END PAR_IN2[8]
  PIN PAR_IN2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 362.885 149.410 366.885 ;
    END
  END PAR_IN2[9]
  PIN PAR_IN3[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 318.960 356.165 319.560 ;
    END
  END PAR_IN3[0]
  PIN PAR_IN3[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END PAR_IN3[10]
  PIN PAR_IN3[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END PAR_IN3[11]
  PIN PAR_IN3[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 362.885 85.930 366.885 ;
    END
  END PAR_IN3[12]
  PIN PAR_IN3[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 113.600 356.165 114.200 ;
    END
  END PAR_IN3[13]
  PIN PAR_IN3[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 178.200 356.165 178.800 ;
    END
  END PAR_IN3[14]
  PIN PAR_IN3[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END PAR_IN3[15]
  PIN PAR_IN3[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 55.120 356.165 55.720 ;
    END
  END PAR_IN3[16]
  PIN PAR_IN3[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 37.440 356.165 38.040 ;
    END
  END PAR_IN3[17]
  PIN PAR_IN3[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END PAR_IN3[18]
  PIN PAR_IN3[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.010 362.885 185.290 366.885 ;
    END
  END PAR_IN3[19]
  PIN PAR_IN3[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.450 362.885 260.730 366.885 ;
    END
  END PAR_IN3[1]
  PIN PAR_IN3[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END PAR_IN3[20]
  PIN PAR_IN3[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END PAR_IN3[21]
  PIN PAR_IN3[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END PAR_IN3[22]
  PIN PAR_IN3[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 289.720 356.165 290.320 ;
    END
  END PAR_IN3[23]
  PIN PAR_IN3[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.510 362.885 288.790 366.885 ;
    END
  END PAR_IN3[24]
  PIN PAR_IN3[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 362.885 117.670 366.885 ;
    END
  END PAR_IN3[25]
  PIN PAR_IN3[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.930 362.885 209.210 366.885 ;
    END
  END PAR_IN3[26]
  PIN PAR_IN3[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END PAR_IN3[27]
  PIN PAR_IN3[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END PAR_IN3[28]
  PIN PAR_IN3[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END PAR_IN3[29]
  PIN PAR_IN3[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 84.360 356.165 84.960 ;
    END
  END PAR_IN3[2]
  PIN PAR_IN3[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 342.760 356.165 343.360 ;
    END
  END PAR_IN3[30]
  PIN PAR_IN3[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 332.210 362.885 332.490 366.885 ;
    END
  END PAR_IN3[31]
  PIN PAR_IN3[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 19.760 356.165 20.360 ;
    END
  END PAR_IN3[3]
  PIN PAR_IN3[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END PAR_IN3[4]
  PIN PAR_IN3[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END PAR_IN3[5]
  PIN PAR_IN3[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END PAR_IN3[6]
  PIN PAR_IN3[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 142.840 356.165 143.440 ;
    END
  END PAR_IN3[7]
  PIN PAR_IN3[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END PAR_IN3[8]
  PIN PAR_IN3[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 360.440 356.165 361.040 ;
    END
  END PAR_IN3[9]
  PIN PAR_IN4[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.850 362.885 233.130 366.885 ;
    END
  END PAR_IN4[0]
  PIN PAR_IN4[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END PAR_IN4[10]
  PIN PAR_IN4[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END PAR_IN4[11]
  PIN PAR_IN4[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 362.885 54.190 366.885 ;
    END
  END PAR_IN4[12]
  PIN PAR_IN4[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END PAR_IN4[13]
  PIN PAR_IN4[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.230 362.885 280.510 366.885 ;
    END
  END PAR_IN4[14]
  PIN PAR_IN4[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END PAR_IN4[15]
  PIN PAR_IN4[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END PAR_IN4[16]
  PIN PAR_IN4[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END PAR_IN4[17]
  PIN PAR_IN4[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END PAR_IN4[18]
  PIN PAR_IN4[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END PAR_IN4[19]
  PIN PAR_IN4[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END PAR_IN4[1]
  PIN PAR_IN4[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.890 362.885 221.170 366.885 ;
    END
  END PAR_IN4[20]
  PIN PAR_IN4[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END PAR_IN4[21]
  PIN PAR_IN4[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.570 362.885 224.850 366.885 ;
    END
  END PAR_IN4[22]
  PIN PAR_IN4[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.110 362.885 316.390 366.885 ;
    END
  END PAR_IN4[23]
  PIN PAR_IN4[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 272.040 356.165 272.640 ;
    END
  END PAR_IN4[24]
  PIN PAR_IN4[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 153.270 362.885 153.550 366.885 ;
    END
  END PAR_IN4[25]
  PIN PAR_IN4[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 155.080 356.165 155.680 ;
    END
  END PAR_IN4[26]
  PIN PAR_IN4[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END PAR_IN4[27]
  PIN PAR_IN4[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END PAR_IN4[28]
  PIN PAR_IN4[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 362.885 2.670 366.885 ;
    END
  END PAR_IN4[29]
  PIN PAR_IN4[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END PAR_IN4[2]
  PIN PAR_IN4[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 13.640 356.165 14.240 ;
    END
  END PAR_IN4[30]
  PIN PAR_IN4[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END PAR_IN4[31]
  PIN PAR_IN4[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.410 362.885 157.690 366.885 ;
    END
  END PAR_IN4[3]
  PIN PAR_IN4[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END PAR_IN4[4]
  PIN PAR_IN4[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 166.640 356.165 167.240 ;
    END
  END PAR_IN4[5]
  PIN PAR_IN4[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END PAR_IN4[6]
  PIN PAR_IN4[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END PAR_IN4[7]
  PIN PAR_IN4[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 362.885 50.050 366.885 ;
    END
  END PAR_IN4[8]
  PIN PAR_IN4[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END PAR_IN4[9]
  PIN PAR_IN5[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END PAR_IN5[0]
  PIN PAR_IN5[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END PAR_IN5[10]
  PIN PAR_IN5[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 66.680 356.165 67.280 ;
    END
  END PAR_IN5[11]
  PIN PAR_IN5[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.530 362.885 236.810 366.885 ;
    END
  END PAR_IN5[12]
  PIN PAR_IN5[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END PAR_IN5[13]
  PIN PAR_IN5[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END PAR_IN5[14]
  PIN PAR_IN5[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END PAR_IN5[15]
  PIN PAR_IN5[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END PAR_IN5[16]
  PIN PAR_IN5[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END PAR_IN5[17]
  PIN PAR_IN5[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.290 362.885 308.570 366.885 ;
    END
  END PAR_IN5[18]
  PIN PAR_IN5[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.110 362.885 201.390 366.885 ;
    END
  END PAR_IN5[19]
  PIN PAR_IN5[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.370 362.885 169.650 366.885 ;
    END
  END PAR_IN5[1]
  PIN PAR_IN5[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 195.880 356.165 196.480 ;
    END
  END PAR_IN5[20]
  PIN PAR_IN5[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.870 362.885 181.150 366.885 ;
    END
  END PAR_IN5[21]
  PIN PAR_IN5[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END PAR_IN5[22]
  PIN PAR_IN5[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 301.280 356.165 301.880 ;
    END
  END PAR_IN5[23]
  PIN PAR_IN5[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 49.000 356.165 49.600 ;
    END
  END PAR_IN5[24]
  PIN PAR_IN5[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END PAR_IN5[25]
  PIN PAR_IN5[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END PAR_IN5[26]
  PIN PAR_IN5[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END PAR_IN5[27]
  PIN PAR_IN5[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END PAR_IN5[28]
  PIN PAR_IN5[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.210 362.885 10.490 366.885 ;
    END
  END PAR_IN5[29]
  PIN PAR_IN5[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 119.720 356.165 120.320 ;
    END
  END PAR_IN5[2]
  PIN PAR_IN5[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END PAR_IN5[30]
  PIN PAR_IN5[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END PAR_IN5[31]
  PIN PAR_IN5[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END PAR_IN5[3]
  PIN PAR_IN5[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.670 362.885 355.950 366.885 ;
    END
  END PAR_IN5[4]
  PIN PAR_IN5[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.190 362.885 292.470 366.885 ;
    END
  END PAR_IN5[5]
  PIN PAR_IN5[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 219.680 356.165 220.280 ;
    END
  END PAR_IN5[6]
  PIN PAR_IN5[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 362.885 137.450 366.885 ;
    END
  END PAR_IN5[7]
  PIN PAR_IN5[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END PAR_IN5[8]
  PIN PAR_IN5[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.810 362.885 245.090 366.885 ;
    END
  END PAR_IN5[9]
  PIN PAR_IN6[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 248.920 356.165 249.520 ;
    END
  END PAR_IN6[0]
  PIN PAR_IN6[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.990 362.885 352.270 366.885 ;
    END
  END PAR_IN6[10]
  PIN PAR_IN6[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 278.160 356.165 278.760 ;
    END
  END PAR_IN6[11]
  PIN PAR_IN6[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 137.400 356.165 138.000 ;
    END
  END PAR_IN6[12]
  PIN PAR_IN6[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 362.885 62.010 366.885 ;
    END
  END PAR_IN6[13]
  PIN PAR_IN6[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 362.885 30.270 366.885 ;
    END
  END PAR_IN6[14]
  PIN PAR_IN6[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 362.885 18.310 366.885 ;
    END
  END PAR_IN6[15]
  PIN PAR_IN6[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END PAR_IN6[16]
  PIN PAR_IN6[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END PAR_IN6[17]
  PIN PAR_IN6[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 307.400 356.165 308.000 ;
    END
  END PAR_IN6[18]
  PIN PAR_IN6[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END PAR_IN6[19]
  PIN PAR_IN6[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END PAR_IN6[1]
  PIN PAR_IN6[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END PAR_IN6[20]
  PIN PAR_IN6[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END PAR_IN6[21]
  PIN PAR_IN6[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 362.885 93.750 366.885 ;
    END
  END PAR_IN6[22]
  PIN PAR_IN6[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.750 362.885 217.030 366.885 ;
    END
  END PAR_IN6[23]
  PIN PAR_IN6[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 354.320 356.165 354.920 ;
    END
  END PAR_IN6[24]
  PIN PAR_IN6[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.890 362.885 336.170 366.885 ;
    END
  END PAR_IN6[25]
  PIN PAR_IN6[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END PAR_IN6[26]
  PIN PAR_IN6[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 295.840 356.165 296.440 ;
    END
  END PAR_IN6[27]
  PIN PAR_IN6[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.550 362.885 276.830 366.885 ;
    END
  END PAR_IN6[28]
  PIN PAR_IN6[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END PAR_IN6[29]
  PIN PAR_IN6[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END PAR_IN6[2]
  PIN PAR_IN6[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END PAR_IN6[30]
  PIN PAR_IN6[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 72.800 356.165 73.400 ;
    END
  END PAR_IN6[31]
  PIN PAR_IN6[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 336.640 356.165 337.240 ;
    END
  END PAR_IN6[3]
  PIN PAR_IN6[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.150 362.885 189.430 366.885 ;
    END
  END PAR_IN6[4]
  PIN PAR_IN6[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 284.280 356.165 284.880 ;
    END
  END PAR_IN6[5]
  PIN PAR_IN6[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END PAR_IN6[6]
  PIN PAR_IN6[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.470 362.885 300.750 366.885 ;
    END
  END PAR_IN6[7]
  PIN PAR_IN6[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.190 362.885 177.470 366.885 ;
    END
  END PAR_IN6[8]
  PIN PAR_IN6[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 313.520 356.165 314.120 ;
    END
  END PAR_IN6[9]
  PIN PAR_IN7[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.170 362.885 344.450 366.885 ;
    END
  END PAR_IN7[0]
  PIN PAR_IN7[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END PAR_IN7[10]
  PIN PAR_IN7[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END PAR_IN7[11]
  PIN PAR_IN7[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END PAR_IN7[12]
  PIN PAR_IN7[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.090 362.885 161.370 366.885 ;
    END
  END PAR_IN7[13]
  PIN PAR_IN7[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END PAR_IN7[14]
  PIN PAR_IN7[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 189.760 356.165 190.360 ;
    END
  END PAR_IN7[15]
  PIN PAR_IN7[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END PAR_IN7[16]
  PIN PAR_IN7[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END PAR_IN7[17]
  PIN PAR_IN7[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END PAR_IN7[18]
  PIN PAR_IN7[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.930 362.885 324.210 366.885 ;
    END
  END PAR_IN7[19]
  PIN PAR_IN7[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 252.630 362.885 252.910 366.885 ;
    END
  END PAR_IN7[1]
  PIN PAR_IN7[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END PAR_IN7[20]
  PIN PAR_IN7[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END PAR_IN7[21]
  PIN PAR_IN7[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.170 362.885 22.450 366.885 ;
    END
  END PAR_IN7[22]
  PIN PAR_IN7[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END PAR_IN7[23]
  PIN PAR_IN7[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END PAR_IN7[24]
  PIN PAR_IN7[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 362.885 296.610 366.885 ;
    END
  END PAR_IN7[25]
  PIN PAR_IN7[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 172.080 356.165 172.680 ;
    END
  END PAR_IN7[26]
  PIN PAR_IN7[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END PAR_IN7[27]
  PIN PAR_IN7[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END PAR_IN7[28]
  PIN PAR_IN7[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 8.200 356.165 8.800 ;
    END
  END PAR_IN7[29]
  PIN PAR_IN7[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END PAR_IN7[2]
  PIN PAR_IN7[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 95.920 356.165 96.520 ;
    END
  END PAR_IN7[30]
  PIN PAR_IN7[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END PAR_IN7[31]
  PIN PAR_IN7[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.150 362.885 304.430 366.885 ;
    END
  END PAR_IN7[3]
  PIN PAR_IN7[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END PAR_IN7[4]
  PIN PAR_IN7[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 184.320 356.165 184.920 ;
    END
  END PAR_IN7[5]
  PIN PAR_IN7[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 362.885 90.070 366.885 ;
    END
  END PAR_IN7[6]
  PIN PAR_IN7[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 362.885 26.590 366.885 ;
    END
  END PAR_IN7[7]
  PIN PAR_IN7[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END PAR_IN7[8]
  PIN PAR_IN7[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.670 362.885 240.950 366.885 ;
    END
  END PAR_IN7[9]
  PIN PAR_IN8[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END PAR_IN8[0]
  PIN PAR_IN8[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 148.960 356.165 149.560 ;
    END
  END PAR_IN8[10]
  PIN PAR_IN8[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END PAR_IN8[11]
  PIN PAR_IN8[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END PAR_IN8[12]
  PIN PAR_IN8[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 362.885 113.990 366.885 ;
    END
  END PAR_IN8[13]
  PIN PAR_IN8[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.230 362.885 165.510 366.885 ;
    END
  END PAR_IN8[14]
  PIN PAR_IN8[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END PAR_IN8[15]
  PIN PAR_IN8[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 348.880 356.165 349.480 ;
    END
  END PAR_IN8[16]
  PIN PAR_IN8[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END PAR_IN8[17]
  PIN PAR_IN8[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END PAR_IN8[18]
  PIN PAR_IN8[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 362.885 38.090 366.885 ;
    END
  END PAR_IN8[19]
  PIN PAR_IN8[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END PAR_IN8[1]
  PIN PAR_IN8[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.970 362.885 312.250 366.885 ;
    END
  END PAR_IN8[20]
  PIN PAR_IN8[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END PAR_IN8[21]
  PIN PAR_IN8[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 225.120 356.165 225.720 ;
    END
  END PAR_IN8[22]
  PIN PAR_IN8[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END PAR_IN8[23]
  PIN PAR_IN8[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 78.240 356.165 78.840 ;
    END
  END PAR_IN8[24]
  PIN PAR_IN8[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END PAR_IN8[25]
  PIN PAR_IN8[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 268.270 362.885 268.550 366.885 ;
    END
  END PAR_IN8[26]
  PIN PAR_IN8[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END PAR_IN8[27]
  PIN PAR_IN8[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 362.885 109.850 366.885 ;
    END
  END PAR_IN8[28]
  PIN PAR_IN8[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END PAR_IN8[29]
  PIN PAR_IN8[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END PAR_IN8[2]
  PIN PAR_IN8[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END PAR_IN8[30]
  PIN PAR_IN8[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 228.710 362.885 228.990 366.885 ;
    END
  END PAR_IN8[31]
  PIN PAR_IN8[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 362.885 70.290 366.885 ;
    END
  END PAR_IN8[3]
  PIN PAR_IN8[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END PAR_IN8[4]
  PIN PAR_IN8[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 362.885 73.970 366.885 ;
    END
  END PAR_IN8[5]
  PIN PAR_IN8[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 107.480 356.165 108.080 ;
    END
  END PAR_IN8[6]
  PIN PAR_IN8[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 90.480 356.165 91.080 ;
    END
  END PAR_IN8[7]
  PIN PAR_IN8[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END PAR_IN8[8]
  PIN PAR_IN8[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.590 362.885 264.870 366.885 ;
    END
  END PAR_IN8[9]
  PIN READY
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.310 362.885 141.590 366.885 ;
    END
  END READY
  PIN RESET
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 362.885 197.250 366.885 ;
    END
  END RESET
  PIN SAMPLE_COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 2.080 356.165 2.680 ;
    END
  END SAMPLE_COUNT[0]
  PIN SAMPLE_COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END SAMPLE_COUNT[1]
  PIN SAMPLE_COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 352.165 266.600 356.165 267.200 ;
    END
  END SAMPLE_COUNT[2]
  PIN SAMPLE_COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END SAMPLE_COUNT[3]
  PIN SERIAL_IN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END SERIAL_IN
  PIN VDD
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 350.520 28.090 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 350.520 104.680 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 5.520 0.085 350.520 353.685 ;
      LAYER met1 ;
        RECT 0.070 0.040 354.590 363.760 ;
      LAYER met2 ;
        RECT 0.090 362.605 2.110 363.790 ;
        RECT 2.950 362.605 5.790 363.790 ;
        RECT 6.630 362.605 9.930 363.790 ;
        RECT 10.770 362.605 14.070 363.790 ;
        RECT 14.910 362.605 17.750 363.790 ;
        RECT 18.590 362.605 21.890 363.790 ;
        RECT 22.730 362.605 26.030 363.790 ;
        RECT 26.870 362.605 29.710 363.790 ;
        RECT 30.550 362.605 33.850 363.790 ;
        RECT 34.690 362.605 37.530 363.790 ;
        RECT 38.370 362.605 41.670 363.790 ;
        RECT 42.510 362.605 45.810 363.790 ;
        RECT 46.650 362.605 49.490 363.790 ;
        RECT 50.330 362.605 53.630 363.790 ;
        RECT 54.470 362.605 57.770 363.790 ;
        RECT 58.610 362.605 61.450 363.790 ;
        RECT 62.290 362.605 65.590 363.790 ;
        RECT 66.430 362.605 69.730 363.790 ;
        RECT 70.570 362.605 73.410 363.790 ;
        RECT 74.250 362.605 77.550 363.790 ;
        RECT 78.390 362.605 81.230 363.790 ;
        RECT 82.070 362.605 85.370 363.790 ;
        RECT 86.210 362.605 89.510 363.790 ;
        RECT 90.350 362.605 93.190 363.790 ;
        RECT 94.030 362.605 97.330 363.790 ;
        RECT 98.170 362.605 101.470 363.790 ;
        RECT 102.310 362.605 105.150 363.790 ;
        RECT 105.990 362.605 109.290 363.790 ;
        RECT 110.130 362.605 113.430 363.790 ;
        RECT 114.270 362.605 117.110 363.790 ;
        RECT 117.950 362.605 121.250 363.790 ;
        RECT 122.090 362.605 124.930 363.790 ;
        RECT 125.770 362.605 129.070 363.790 ;
        RECT 129.910 362.605 133.210 363.790 ;
        RECT 134.050 362.605 136.890 363.790 ;
        RECT 137.730 362.605 141.030 363.790 ;
        RECT 141.870 362.605 145.170 363.790 ;
        RECT 146.010 362.605 148.850 363.790 ;
        RECT 149.690 362.605 152.990 363.790 ;
        RECT 153.830 362.605 157.130 363.790 ;
        RECT 157.970 362.605 160.810 363.790 ;
        RECT 161.650 362.605 164.950 363.790 ;
        RECT 165.790 362.605 169.090 363.790 ;
        RECT 169.930 362.605 172.770 363.790 ;
        RECT 173.610 362.605 176.910 363.790 ;
        RECT 177.750 362.605 180.590 363.790 ;
        RECT 181.430 362.605 184.730 363.790 ;
        RECT 185.570 362.605 188.870 363.790 ;
        RECT 189.710 362.605 192.550 363.790 ;
        RECT 193.390 362.605 196.690 363.790 ;
        RECT 197.530 362.605 200.830 363.790 ;
        RECT 201.670 362.605 204.510 363.790 ;
        RECT 205.350 362.605 208.650 363.790 ;
        RECT 209.490 362.605 212.790 363.790 ;
        RECT 213.630 362.605 216.470 363.790 ;
        RECT 217.310 362.605 220.610 363.790 ;
        RECT 221.450 362.605 224.290 363.790 ;
        RECT 225.130 362.605 228.430 363.790 ;
        RECT 229.270 362.605 232.570 363.790 ;
        RECT 233.410 362.605 236.250 363.790 ;
        RECT 237.090 362.605 240.390 363.790 ;
        RECT 241.230 362.605 244.530 363.790 ;
        RECT 245.370 362.605 248.210 363.790 ;
        RECT 249.050 362.605 252.350 363.790 ;
        RECT 253.190 362.605 256.490 363.790 ;
        RECT 257.330 362.605 260.170 363.790 ;
        RECT 261.010 362.605 264.310 363.790 ;
        RECT 265.150 362.605 267.990 363.790 ;
        RECT 268.830 362.605 272.130 363.790 ;
        RECT 272.970 362.605 276.270 363.790 ;
        RECT 277.110 362.605 279.950 363.790 ;
        RECT 280.790 362.605 284.090 363.790 ;
        RECT 284.930 362.605 288.230 363.790 ;
        RECT 289.070 362.605 291.910 363.790 ;
        RECT 292.750 362.605 296.050 363.790 ;
        RECT 296.890 362.605 300.190 363.790 ;
        RECT 301.030 362.605 303.870 363.790 ;
        RECT 304.710 362.605 308.010 363.790 ;
        RECT 308.850 362.605 311.690 363.790 ;
        RECT 312.530 362.605 315.830 363.790 ;
        RECT 316.670 362.605 319.970 363.790 ;
        RECT 320.810 362.605 323.650 363.790 ;
        RECT 324.490 362.605 327.790 363.790 ;
        RECT 328.630 362.605 331.930 363.790 ;
        RECT 332.770 362.605 335.610 363.790 ;
        RECT 336.450 362.605 339.750 363.790 ;
        RECT 340.590 362.605 343.890 363.790 ;
        RECT 344.730 362.605 347.570 363.790 ;
        RECT 348.410 362.605 351.710 363.790 ;
        RECT 352.550 362.605 355.390 363.790 ;
        RECT 0.090 4.280 355.670 362.605 ;
        RECT 0.650 0.010 3.490 4.280 ;
        RECT 4.330 0.010 7.630 4.280 ;
        RECT 8.470 0.010 11.310 4.280 ;
        RECT 12.150 0.010 15.450 4.280 ;
        RECT 16.290 0.010 19.590 4.280 ;
        RECT 20.430 0.010 23.270 4.280 ;
        RECT 24.110 0.010 27.410 4.280 ;
        RECT 28.250 0.010 31.550 4.280 ;
        RECT 32.390 0.010 35.230 4.280 ;
        RECT 36.070 0.010 39.370 4.280 ;
        RECT 40.210 0.010 43.510 4.280 ;
        RECT 44.350 0.010 47.190 4.280 ;
        RECT 48.030 0.010 51.330 4.280 ;
        RECT 52.170 0.010 55.010 4.280 ;
        RECT 55.850 0.010 59.150 4.280 ;
        RECT 59.990 0.010 63.290 4.280 ;
        RECT 64.130 0.010 66.970 4.280 ;
        RECT 67.810 0.010 71.110 4.280 ;
        RECT 71.950 0.010 75.250 4.280 ;
        RECT 76.090 0.010 78.930 4.280 ;
        RECT 79.770 0.010 83.070 4.280 ;
        RECT 83.910 0.010 87.210 4.280 ;
        RECT 88.050 0.010 90.890 4.280 ;
        RECT 91.730 0.010 95.030 4.280 ;
        RECT 95.870 0.010 98.710 4.280 ;
        RECT 99.550 0.010 102.850 4.280 ;
        RECT 103.690 0.010 106.990 4.280 ;
        RECT 107.830 0.010 110.670 4.280 ;
        RECT 111.510 0.010 114.810 4.280 ;
        RECT 115.650 0.010 118.950 4.280 ;
        RECT 119.790 0.010 122.630 4.280 ;
        RECT 123.470 0.010 126.770 4.280 ;
        RECT 127.610 0.010 130.910 4.280 ;
        RECT 131.750 0.010 134.590 4.280 ;
        RECT 135.430 0.010 138.730 4.280 ;
        RECT 139.570 0.010 142.410 4.280 ;
        RECT 143.250 0.010 146.550 4.280 ;
        RECT 147.390 0.010 150.690 4.280 ;
        RECT 151.530 0.010 154.370 4.280 ;
        RECT 155.210 0.010 158.510 4.280 ;
        RECT 159.350 0.010 162.650 4.280 ;
        RECT 163.490 0.010 166.330 4.280 ;
        RECT 167.170 0.010 170.470 4.280 ;
        RECT 171.310 0.010 174.610 4.280 ;
        RECT 175.450 0.010 178.290 4.280 ;
        RECT 179.130 0.010 182.430 4.280 ;
        RECT 183.270 0.010 186.110 4.280 ;
        RECT 186.950 0.010 190.250 4.280 ;
        RECT 191.090 0.010 194.390 4.280 ;
        RECT 195.230 0.010 198.070 4.280 ;
        RECT 198.910 0.010 202.210 4.280 ;
        RECT 203.050 0.010 206.350 4.280 ;
        RECT 207.190 0.010 210.030 4.280 ;
        RECT 210.870 0.010 214.170 4.280 ;
        RECT 215.010 0.010 218.310 4.280 ;
        RECT 219.150 0.010 221.990 4.280 ;
        RECT 222.830 0.010 226.130 4.280 ;
        RECT 226.970 0.010 230.270 4.280 ;
        RECT 231.110 0.010 233.950 4.280 ;
        RECT 234.790 0.010 238.090 4.280 ;
        RECT 238.930 0.010 241.770 4.280 ;
        RECT 242.610 0.010 245.910 4.280 ;
        RECT 246.750 0.010 250.050 4.280 ;
        RECT 250.890 0.010 253.730 4.280 ;
        RECT 254.570 0.010 257.870 4.280 ;
        RECT 258.710 0.010 262.010 4.280 ;
        RECT 262.850 0.010 265.690 4.280 ;
        RECT 266.530 0.010 269.830 4.280 ;
        RECT 270.670 0.010 273.970 4.280 ;
        RECT 274.810 0.010 277.650 4.280 ;
        RECT 278.490 0.010 281.790 4.280 ;
        RECT 282.630 0.010 285.470 4.280 ;
        RECT 286.310 0.010 289.610 4.280 ;
        RECT 290.450 0.010 293.750 4.280 ;
        RECT 294.590 0.010 297.430 4.280 ;
        RECT 298.270 0.010 301.570 4.280 ;
        RECT 302.410 0.010 305.710 4.280 ;
        RECT 306.550 0.010 309.390 4.280 ;
        RECT 310.230 0.010 313.530 4.280 ;
        RECT 314.370 0.010 317.670 4.280 ;
        RECT 318.510 0.010 321.350 4.280 ;
        RECT 322.190 0.010 325.490 4.280 ;
        RECT 326.330 0.010 329.170 4.280 ;
        RECT 330.010 0.010 333.310 4.280 ;
        RECT 334.150 0.010 337.450 4.280 ;
        RECT 338.290 0.010 341.130 4.280 ;
        RECT 341.970 0.010 345.270 4.280 ;
        RECT 346.110 0.010 349.410 4.280 ;
        RECT 350.250 0.010 353.090 4.280 ;
        RECT 353.930 0.010 355.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 363.440 353.010 363.840 ;
        RECT 0.310 361.440 353.010 363.440 ;
        RECT 0.310 360.040 351.765 361.440 ;
        RECT 0.310 358.720 353.010 360.040 ;
        RECT 4.400 357.320 353.010 358.720 ;
        RECT 0.310 355.320 353.010 357.320 ;
        RECT 0.310 353.920 351.765 355.320 ;
        RECT 0.310 353.280 353.010 353.920 ;
        RECT 4.400 351.880 353.010 353.280 ;
        RECT 0.310 349.880 353.010 351.880 ;
        RECT 0.310 348.480 351.765 349.880 ;
        RECT 0.310 347.160 353.010 348.480 ;
        RECT 4.400 345.760 353.010 347.160 ;
        RECT 0.310 343.760 353.010 345.760 ;
        RECT 0.310 342.360 351.765 343.760 ;
        RECT 0.310 341.720 353.010 342.360 ;
        RECT 4.400 340.320 353.010 341.720 ;
        RECT 0.310 337.640 353.010 340.320 ;
        RECT 0.310 336.240 351.765 337.640 ;
        RECT 0.310 335.600 353.010 336.240 ;
        RECT 4.400 334.200 353.010 335.600 ;
        RECT 0.310 332.200 353.010 334.200 ;
        RECT 0.310 330.800 351.765 332.200 ;
        RECT 0.310 329.480 353.010 330.800 ;
        RECT 4.400 328.080 353.010 329.480 ;
        RECT 0.310 326.080 353.010 328.080 ;
        RECT 0.310 324.680 351.765 326.080 ;
        RECT 0.310 324.040 353.010 324.680 ;
        RECT 4.400 322.640 353.010 324.040 ;
        RECT 0.310 319.960 353.010 322.640 ;
        RECT 0.310 318.560 351.765 319.960 ;
        RECT 0.310 317.920 353.010 318.560 ;
        RECT 4.400 316.520 353.010 317.920 ;
        RECT 0.310 314.520 353.010 316.520 ;
        RECT 0.310 313.120 351.765 314.520 ;
        RECT 0.310 311.800 353.010 313.120 ;
        RECT 4.400 310.400 353.010 311.800 ;
        RECT 0.310 308.400 353.010 310.400 ;
        RECT 0.310 307.000 351.765 308.400 ;
        RECT 0.310 306.360 353.010 307.000 ;
        RECT 4.400 304.960 353.010 306.360 ;
        RECT 0.310 302.280 353.010 304.960 ;
        RECT 0.310 300.880 351.765 302.280 ;
        RECT 0.310 300.240 353.010 300.880 ;
        RECT 4.400 298.840 353.010 300.240 ;
        RECT 0.310 296.840 353.010 298.840 ;
        RECT 0.310 295.440 351.765 296.840 ;
        RECT 0.310 294.120 353.010 295.440 ;
        RECT 4.400 292.720 353.010 294.120 ;
        RECT 0.310 290.720 353.010 292.720 ;
        RECT 0.310 289.320 351.765 290.720 ;
        RECT 0.310 288.680 353.010 289.320 ;
        RECT 4.400 287.280 353.010 288.680 ;
        RECT 0.310 285.280 353.010 287.280 ;
        RECT 0.310 283.880 351.765 285.280 ;
        RECT 0.310 282.560 353.010 283.880 ;
        RECT 4.400 281.160 353.010 282.560 ;
        RECT 0.310 279.160 353.010 281.160 ;
        RECT 0.310 277.760 351.765 279.160 ;
        RECT 0.310 276.440 353.010 277.760 ;
        RECT 4.400 275.040 353.010 276.440 ;
        RECT 0.310 273.040 353.010 275.040 ;
        RECT 0.310 271.640 351.765 273.040 ;
        RECT 0.310 271.000 353.010 271.640 ;
        RECT 4.400 269.600 353.010 271.000 ;
        RECT 0.310 267.600 353.010 269.600 ;
        RECT 0.310 266.200 351.765 267.600 ;
        RECT 0.310 264.880 353.010 266.200 ;
        RECT 4.400 263.480 353.010 264.880 ;
        RECT 0.310 261.480 353.010 263.480 ;
        RECT 0.310 260.080 351.765 261.480 ;
        RECT 0.310 259.440 353.010 260.080 ;
        RECT 4.400 258.040 353.010 259.440 ;
        RECT 0.310 255.360 353.010 258.040 ;
        RECT 0.310 253.960 351.765 255.360 ;
        RECT 0.310 253.320 353.010 253.960 ;
        RECT 4.400 251.920 353.010 253.320 ;
        RECT 0.310 249.920 353.010 251.920 ;
        RECT 0.310 248.520 351.765 249.920 ;
        RECT 0.310 247.200 353.010 248.520 ;
        RECT 4.400 245.800 353.010 247.200 ;
        RECT 0.310 243.800 353.010 245.800 ;
        RECT 0.310 242.400 351.765 243.800 ;
        RECT 0.310 241.760 353.010 242.400 ;
        RECT 4.400 240.360 353.010 241.760 ;
        RECT 0.310 237.680 353.010 240.360 ;
        RECT 0.310 236.280 351.765 237.680 ;
        RECT 0.310 235.640 353.010 236.280 ;
        RECT 4.400 234.240 353.010 235.640 ;
        RECT 0.310 232.240 353.010 234.240 ;
        RECT 0.310 230.840 351.765 232.240 ;
        RECT 0.310 229.520 353.010 230.840 ;
        RECT 4.400 228.120 353.010 229.520 ;
        RECT 0.310 226.120 353.010 228.120 ;
        RECT 0.310 224.720 351.765 226.120 ;
        RECT 0.310 224.080 353.010 224.720 ;
        RECT 4.400 222.680 353.010 224.080 ;
        RECT 0.310 220.680 353.010 222.680 ;
        RECT 0.310 219.280 351.765 220.680 ;
        RECT 0.310 217.960 353.010 219.280 ;
        RECT 4.400 216.560 353.010 217.960 ;
        RECT 0.310 214.560 353.010 216.560 ;
        RECT 0.310 213.160 351.765 214.560 ;
        RECT 0.310 211.840 353.010 213.160 ;
        RECT 4.400 210.440 353.010 211.840 ;
        RECT 0.310 208.440 353.010 210.440 ;
        RECT 0.310 207.040 351.765 208.440 ;
        RECT 0.310 206.400 353.010 207.040 ;
        RECT 4.400 205.000 353.010 206.400 ;
        RECT 0.310 203.000 353.010 205.000 ;
        RECT 0.310 201.600 351.765 203.000 ;
        RECT 0.310 200.280 353.010 201.600 ;
        RECT 4.400 198.880 353.010 200.280 ;
        RECT 0.310 196.880 353.010 198.880 ;
        RECT 0.310 195.480 351.765 196.880 ;
        RECT 0.310 194.840 353.010 195.480 ;
        RECT 4.400 193.440 353.010 194.840 ;
        RECT 0.310 190.760 353.010 193.440 ;
        RECT 0.310 189.360 351.765 190.760 ;
        RECT 0.310 188.720 353.010 189.360 ;
        RECT 4.400 187.320 353.010 188.720 ;
        RECT 0.310 185.320 353.010 187.320 ;
        RECT 0.310 183.920 351.765 185.320 ;
        RECT 0.310 182.600 353.010 183.920 ;
        RECT 4.400 181.200 353.010 182.600 ;
        RECT 0.310 179.200 353.010 181.200 ;
        RECT 0.310 177.800 351.765 179.200 ;
        RECT 0.310 177.160 353.010 177.800 ;
        RECT 4.400 175.760 353.010 177.160 ;
        RECT 0.310 173.080 353.010 175.760 ;
        RECT 0.310 171.680 351.765 173.080 ;
        RECT 0.310 171.040 353.010 171.680 ;
        RECT 4.400 169.640 353.010 171.040 ;
        RECT 0.310 167.640 353.010 169.640 ;
        RECT 0.310 166.240 351.765 167.640 ;
        RECT 0.310 164.920 353.010 166.240 ;
        RECT 4.400 163.520 353.010 164.920 ;
        RECT 0.310 161.520 353.010 163.520 ;
        RECT 0.310 160.120 351.765 161.520 ;
        RECT 0.310 159.480 353.010 160.120 ;
        RECT 4.400 158.080 353.010 159.480 ;
        RECT 0.310 156.080 353.010 158.080 ;
        RECT 0.310 154.680 351.765 156.080 ;
        RECT 0.310 153.360 353.010 154.680 ;
        RECT 4.400 151.960 353.010 153.360 ;
        RECT 0.310 149.960 353.010 151.960 ;
        RECT 0.310 148.560 351.765 149.960 ;
        RECT 0.310 147.240 353.010 148.560 ;
        RECT 4.400 145.840 353.010 147.240 ;
        RECT 0.310 143.840 353.010 145.840 ;
        RECT 0.310 142.440 351.765 143.840 ;
        RECT 0.310 141.800 353.010 142.440 ;
        RECT 4.400 140.400 353.010 141.800 ;
        RECT 0.310 138.400 353.010 140.400 ;
        RECT 0.310 137.000 351.765 138.400 ;
        RECT 0.310 135.680 353.010 137.000 ;
        RECT 4.400 134.280 353.010 135.680 ;
        RECT 0.310 132.280 353.010 134.280 ;
        RECT 0.310 130.880 351.765 132.280 ;
        RECT 0.310 130.240 353.010 130.880 ;
        RECT 4.400 128.840 353.010 130.240 ;
        RECT 0.310 126.160 353.010 128.840 ;
        RECT 0.310 124.760 351.765 126.160 ;
        RECT 0.310 124.120 353.010 124.760 ;
        RECT 4.400 122.720 353.010 124.120 ;
        RECT 0.310 120.720 353.010 122.720 ;
        RECT 0.310 119.320 351.765 120.720 ;
        RECT 0.310 118.000 353.010 119.320 ;
        RECT 4.400 116.600 353.010 118.000 ;
        RECT 0.310 114.600 353.010 116.600 ;
        RECT 0.310 113.200 351.765 114.600 ;
        RECT 0.310 112.560 353.010 113.200 ;
        RECT 4.400 111.160 353.010 112.560 ;
        RECT 0.310 108.480 353.010 111.160 ;
        RECT 0.310 107.080 351.765 108.480 ;
        RECT 0.310 106.440 353.010 107.080 ;
        RECT 4.400 105.040 353.010 106.440 ;
        RECT 0.310 103.040 353.010 105.040 ;
        RECT 0.310 101.640 351.765 103.040 ;
        RECT 0.310 100.320 353.010 101.640 ;
        RECT 4.400 98.920 353.010 100.320 ;
        RECT 0.310 96.920 353.010 98.920 ;
        RECT 0.310 95.520 351.765 96.920 ;
        RECT 0.310 94.880 353.010 95.520 ;
        RECT 4.400 93.480 353.010 94.880 ;
        RECT 0.310 91.480 353.010 93.480 ;
        RECT 0.310 90.080 351.765 91.480 ;
        RECT 0.310 88.760 353.010 90.080 ;
        RECT 4.400 87.360 353.010 88.760 ;
        RECT 0.310 85.360 353.010 87.360 ;
        RECT 0.310 83.960 351.765 85.360 ;
        RECT 0.310 82.640 353.010 83.960 ;
        RECT 4.400 81.240 353.010 82.640 ;
        RECT 0.310 79.240 353.010 81.240 ;
        RECT 0.310 77.840 351.765 79.240 ;
        RECT 0.310 77.200 353.010 77.840 ;
        RECT 4.400 75.800 353.010 77.200 ;
        RECT 0.310 73.800 353.010 75.800 ;
        RECT 0.310 72.400 351.765 73.800 ;
        RECT 0.310 71.080 353.010 72.400 ;
        RECT 4.400 69.680 353.010 71.080 ;
        RECT 0.310 67.680 353.010 69.680 ;
        RECT 0.310 66.280 351.765 67.680 ;
        RECT 0.310 65.640 353.010 66.280 ;
        RECT 4.400 64.240 353.010 65.640 ;
        RECT 0.310 61.560 353.010 64.240 ;
        RECT 0.310 60.160 351.765 61.560 ;
        RECT 0.310 59.520 353.010 60.160 ;
        RECT 4.400 58.120 353.010 59.520 ;
        RECT 0.310 56.120 353.010 58.120 ;
        RECT 0.310 54.720 351.765 56.120 ;
        RECT 0.310 53.400 353.010 54.720 ;
        RECT 4.400 52.000 353.010 53.400 ;
        RECT 0.310 50.000 353.010 52.000 ;
        RECT 0.310 48.600 351.765 50.000 ;
        RECT 0.310 47.960 353.010 48.600 ;
        RECT 4.400 46.560 353.010 47.960 ;
        RECT 0.310 43.880 353.010 46.560 ;
        RECT 0.310 42.480 351.765 43.880 ;
        RECT 0.310 41.840 353.010 42.480 ;
        RECT 4.400 40.440 353.010 41.840 ;
        RECT 0.310 38.440 353.010 40.440 ;
        RECT 0.310 37.040 351.765 38.440 ;
        RECT 0.310 35.720 353.010 37.040 ;
        RECT 4.400 34.320 353.010 35.720 ;
        RECT 0.310 32.320 353.010 34.320 ;
        RECT 0.310 30.920 351.765 32.320 ;
        RECT 0.310 30.280 353.010 30.920 ;
        RECT 4.400 28.880 353.010 30.280 ;
        RECT 0.310 26.200 353.010 28.880 ;
        RECT 0.310 24.800 351.765 26.200 ;
        RECT 0.310 24.160 353.010 24.800 ;
        RECT 4.400 22.760 353.010 24.160 ;
        RECT 0.310 20.760 353.010 22.760 ;
        RECT 0.310 19.360 351.765 20.760 ;
        RECT 0.310 18.040 353.010 19.360 ;
        RECT 4.400 16.640 353.010 18.040 ;
        RECT 0.310 14.640 353.010 16.640 ;
        RECT 0.310 13.240 351.765 14.640 ;
        RECT 0.310 12.600 353.010 13.240 ;
        RECT 4.400 11.200 353.010 12.600 ;
        RECT 0.310 9.200 353.010 11.200 ;
        RECT 0.310 7.800 351.765 9.200 ;
        RECT 0.310 6.480 353.010 7.800 ;
        RECT 4.400 5.080 353.010 6.480 ;
        RECT 0.310 3.080 353.010 5.080 ;
        RECT 0.310 2.230 351.765 3.080 ;
      LAYER met4 ;
        RECT 21.040 10.640 352.985 353.840 ;
      LAYER met5 ;
        RECT 5.520 157.300 350.520 334.450 ;
  END
END deserialiser_unit_cell_1
END LIBRARY

