* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599419937836
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_599419937837
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT DFL1sd_CDNS_599419937832
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFL1sd2_CDNS_599419937833
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT Inverter2 GND VDD INP OUT
** N=4 EP=4 IP=31 FDC=28
M0 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=-445 $Y=-6375 $D=9
M1 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=-15 $Y=-6375 $D=9
M2 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=415 $Y=-6375 $D=9
M3 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=845 $Y=-6375 $D=9
M4 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1275 $Y=-6375 $D=9
M5 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1705 $Y=-6375 $D=9
M6 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2135 $Y=-6375 $D=9
M7 GND INP OUT GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2565 $Y=-6375 $D=9
M8 OUT INP GND GND nshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2995 $Y=-6375 $D=9
M9 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=-670 $Y=-110 $D=79
M10 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=-240 $Y=-110 $D=79
M11 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=190 $Y=-110 $D=79
M12 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=620 $Y=-110 $D=79
M13 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1050 $Y=-110 $D=79
M14 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1480 $Y=-110 $D=79
M15 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=1910 $Y=-110 $D=79
M16 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2340 $Y=-110 $D=79
M17 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=2770 $Y=-110 $D=79
M18 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3200 $Y=-110 $D=79
M19 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=3630 $Y=-110 $D=79
M20 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4060 $Y=-110 $D=79
M21 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4490 $Y=-110 $D=79
M22 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=4920 $Y=-110 $D=79
M23 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5350 $Y=-110 $D=79
M24 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=5780 $Y=-110 $D=79
M25 OUT INP VDD VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6210 $Y=-110 $D=79
M26 VDD INP OUT VDD pshort L=0.15 W=5 m=1 r=33.3333 a=0.75 p=10.3 mult=1 $X=6640 $Y=-110 $D=79
X27 GND VDD Dpar a=48.4008 p=28.78 m=1 $[nwdiode] $X=-1795 $Y=-290 $D=185
.ENDS
***************************************
