* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT mrdn POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdn_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp POS NEG SUB
.ENDS
***************************************
.SUBCKT mrdp_hv POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xpwres POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_3 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=0.59 W=0.55 m=1 r=0.932203 a=0.3245 p=2.28 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=0.59 W=0.87 m=1 r=1.47458 a=0.5133 p=2.92 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 1 0 $X=-190 $Y=-2960
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_8 VNB VPB VGND VPWR
** N=16 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=2.89 W=0.55 m=1 r=0.190311 a=1.5895 p=6.88 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=2.89 W=0.87 m=1 r=0.301038 a=2.5143 p=7.52 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_12 VNB VPB VGND VPWR
** N=18 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=4.73 W=0.55 m=1 r=0.116279 a=2.6015 p=10.56 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=4.73 W=0.87 m=1 r=0.183932 a=4.1151 p=11.2 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
** N=12 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.05 W=0.55 m=1 r=0.52381 a=0.5775 p=3.2 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.05 W=0.87 m=1 r=0.828571 a=0.9135 p=3.84 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__diode_2 VNB DIODE
** N=9 EP=2 IP=0 FDC=1
*.SEEDPROM
D0 VNB DIODE ndiode AREA=0.4347 PJ=2.64 m=1 ahftempperim=2.64 $X=155 $Y=195 $D=167
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_6 VNB VPB VGND VPWR
** N=14 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.97 W=0.55 m=1 r=0.279188 a=1.0835 p=5.04 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.97 W=0.87 m=1 r=0.441624 a=1.7139 p=5.68 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_7 1 3 4
** N=4 EP=3 IP=10 FDC=2
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 4 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dfrtp_4 VNB VPB CLK D RESET_B VPWR Q VGND
** N=88 EP=8 IP=0 FDC=34
*.SEEDPROM
M0 VGND CLK 9 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 10 9 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 15 D VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2090 $Y=235 $D=9
M3 12 9 15 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=2565 $Y=235 $D=9
M4 18 10 12 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=3045 $Y=235 $D=9
M5 19 11 18 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3875 $Y=235 $D=8
M6 VGND RESET_B 19 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4235 $Y=235 $D=9
M7 11 12 VGND VNB nshort L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=4895 $Y=235 $D=9
M8 14 10 11 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5390 $Y=235 $D=9
M9 20 9 14 VNB nshort L=0.15 W=0.36 m=1 r=2.4 a=0.054 p=1.02 mult=1 $X=5935 $Y=235 $D=9
M10 VGND 13 20 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M11 21 RESET_B VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=235 $D=9
M12 13 14 21 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7615 $Y=235 $D=9
M13 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8555 $Y=235 $D=9
M14 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=8975 $Y=235 $D=9
M15 Q 13 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9395 $Y=235 $D=9
M16 VGND 13 Q VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=9815 $Y=235 $D=9
M17 VPWR CLK 9 VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M18 10 9 VPWR VPB phighvt L=0.15 W=0.64 m=1 r=4.26667 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M19 15 D VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2150 $Y=2065 $D=89
M20 12 10 15 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2610 $Y=2065 $D=89
M21 16 9 12 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3105 $Y=2065 $D=89
M22 VPWR 11 16 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3805 $Y=2065 $D=89
M23 16 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4290 $Y=2065 $D=89
M24 11 12 VPWR VPB phighvt L=0.15 W=0.84 m=1 r=5.6 a=0.126 p=1.98 mult=1 $X=5275 $Y=1645 $D=89
M25 14 9 11 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5770 $Y=2065 $D=89
M26 17 10 14 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6200 $Y=2065 $D=89
M27 VPWR 13 17 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6620 $Y=2065 $D=89
M28 13 RESET_B VPWR VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7160 $Y=2065 $D=89
M29 VPWR 14 13 VPB phighvt L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7580 $Y=2065 $D=89
M30 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8555 $Y=1485 $D=89
M31 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8975 $Y=1485 $D=89
M32 Q 13 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9395 $Y=1485 $D=89
M33 VPWR 13 Q VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=9815 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_9 $T=5980 0 0 0 $X=5790 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=36
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=10580 0 0 0 $X=10390 $Y=-240
X1 1 2 3 4 6 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_14 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_15 1 3
** N=3 EP=2 IP=7 FDC=1
*.SEEDPROM
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=920 0 0 0 $X=730 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__inv_8 VNB VPB A VPWR Y VGND
** N=48 EP=6 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=560 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=980 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1400 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1820 $Y=235 $D=9
M4 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2240 $Y=235 $D=9
M5 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2660 $Y=235 $D=9
M6 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3080 $Y=235 $D=9
M7 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3500 $Y=235 $D=9
M8 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=560 $Y=1485 $D=89
M9 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=980 $Y=1485 $D=89
M10 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1400 $Y=1485 $D=89
M11 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1820 $Y=1485 $D=89
M12 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2240 $Y=1485 $D=89
M13 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2660 $Y=1485 $D=89
M14 Y A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3080 $Y=1485 $D=89
M15 VPWR A Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3500 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7
** N=7 EP=7 IP=13 FDC=35
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 5 7 2 6 1 sky130_fd_sc_hd__dfrtp_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=34
*.SEEDPROM
X1 1 2 3 4 6 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor2_4 VNB VPB A B VPWR Y VGND
** N=51 EP=7 IP=0 FDC=16
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M9 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M10 VPWR A 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M11 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M12 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M13 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M14 Y B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M15 8 B Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=4 FDC=12
*.SEEDPROM
X0 1 2 ICV_10 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_10 $T=14260 0 0 0 $X=14070 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o22a_4 VNB VPB B1 B2 A1 A2 VPWR X VGND
** N=65 EP=9 IP=0 FDC=24
*.SEEDPROM
M0 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=480 $Y=235 $D=9
M1 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=900 $Y=235 $D=9
M2 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=9
M3 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1740 $Y=235 $D=9
M4 10 B1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2680 $Y=235 $D=9
M5 13 B2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3100 $Y=235 $D=9
M6 10 B2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3520 $Y=235 $D=9
M7 13 B1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3940 $Y=235 $D=9
M8 VGND A1 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4440 $Y=235 $D=9
M9 13 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4860 $Y=235 $D=9
M10 VGND A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5280 $Y=235 $D=9
M11 13 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5700 $Y=235 $D=9
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=480 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=900 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M16 11 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2680 $Y=1485 $D=89
M17 10 B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3100 $Y=1485 $D=89
M18 11 B2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3520 $Y=1485 $D=89
M19 VPWR B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3940 $Y=1485 $D=89
M20 12 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4440 $Y=1485 $D=89
M21 10 A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4860 $Y=1485 $D=89
M22 12 A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5280 $Y=1485 $D=89
M23 VPWR A1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5700 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__buf_1 VNB VPB A VPWR X VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND A 7 VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 X 7 VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR A 7 VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 X 7 VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__o21a_4 VNB VPB B1 A1 A2 VPWR X VGND
** N=53 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 9 B1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2640 $Y=235 $D=9
M5 12 B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3070 $Y=235 $D=9
M6 VGND A1 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M7 12 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4090 $Y=235 $D=9
M8 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4520 $Y=235 $D=9
M9 12 A1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4950 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=720 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1150 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1580 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2010 $Y=1485 $D=89
M14 9 B1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2460 $Y=1485 $D=89
M15 VPWR B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2890 $Y=1485 $D=89
M16 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3660 $Y=1485 $D=89
M17 9 A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4090 $Y=1485 $D=89
M18 11 A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4520 $Y=1485 $D=89
M19 VPWR A1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4950 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251
** N=419 EP=251 IP=4594 FDC=8221
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=314105 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=319545 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=324985 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=330425 $D=191
X4 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=335865 $D=191
X5 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=341305 $D=191
X6 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=346745 $D=191
X7 1 2 Dpar a=554.335 p=693.97 m=1 $[nwdiode] $X=5330 $Y=352185 $D=191
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 340000 0 0 $X=6710 $Y=339760
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 340000 1 0 $X=25570 $Y=337040
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28520 312800 0 0 $X=28330 $Y=312560
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=30360 345440 0 0 $X=30170 $Y=345200
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=32200 329120 0 0 $X=32010 $Y=328880
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=34040 318240 0 0 $X=33850 $Y=318000
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=51980 323680 1 0 $X=51790 $Y=320720
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=54740 340000 0 0 $X=54550 $Y=339760
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=58420 345440 0 0 $X=58230 $Y=345200
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=62100 334560 0 0 $X=61910 $Y=334320
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=72680 340000 1 0 $X=72490 $Y=337040
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74520 312800 1 0 $X=74330 $Y=309840
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74520 334560 1 0 $X=74330 $Y=331600
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74980 345440 0 0 $X=74790 $Y=345200
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=84640 323680 0 0 $X=84450 $Y=323440
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=84640 340000 0 0 $X=84450 $Y=339760
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=86480 318240 0 0 $X=86290 $Y=318000
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=86480 345440 0 0 $X=86290 $Y=345200
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88780 340000 1 0 $X=88590 $Y=337040
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 340000 1 0 $X=102390 $Y=337040
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=108100 345440 1 0 $X=107910 $Y=342480
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=109940 318240 0 0 $X=109750 $Y=318000
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=117300 323680 1 0 $X=117110 $Y=320720
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=121440 334560 1 0 $X=121250 $Y=331600
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=123740 334560 0 0 $X=123550 $Y=334320
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 318240 1 0 $X=130450 $Y=315280
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 350880 1 0 $X=130450 $Y=347920
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=140760 345440 0 0 $X=140570 $Y=345200
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 318240 0 0 $X=144250 $Y=318000
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=146280 329120 1 0 $X=146090 $Y=326160
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=146280 329120 0 0 $X=146090 $Y=328880
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=149960 312800 0 0 $X=149770 $Y=312560
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=155480 312800 1 0 $X=155290 $Y=309840
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=155480 318240 1 0 $X=155290 $Y=315280
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164220 329120 1 0 $X=164030 $Y=326160
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=166060 345440 1 0 $X=165870 $Y=342480
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=166980 318240 0 0 $X=166790 $Y=318000
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=166980 345440 0 0 $X=166790 $Y=345200
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 312800 1 0 $X=174150 $Y=309840
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=182620 329120 1 0 $X=182430 $Y=326160
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=184460 312800 1 0 $X=184270 $Y=309840
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=188600 329120 0 0 $X=188410 $Y=328880
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=188600 334560 1 0 $X=188410 $Y=331600
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=192740 329120 0 0 $X=192550 $Y=328880
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=198720 323680 1 0 $X=198530 $Y=320720
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=200560 334560 0 0 $X=200370 $Y=334320
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=203320 318240 1 0 $X=203130 $Y=315280
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=208840 345440 1 0 $X=208650 $Y=342480
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=211600 334560 1 0 $X=211410 $Y=331600
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 345440 1 0 $X=214630 $Y=342480
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 350880 1 0 $X=214630 $Y=347920
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=216660 312800 1 0 $X=216470 $Y=309840
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=226780 318240 0 0 $X=226590 $Y=318000
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 312800 0 0 $X=230270 $Y=312560
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 323680 1 0 $X=242690 $Y=320720
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 340000 1 0 $X=242690 $Y=337040
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=247020 323680 0 0 $X=246830 $Y=323440
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=250240 340000 1 0 $X=250050 $Y=337040
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=267720 340000 1 0 $X=267530 $Y=337040
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 318240 1 0 $X=270750 $Y=315280
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 323680 1 0 $X=270750 $Y=320720
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=272780 318240 1 0 $X=272590 $Y=315280
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 323680 0 0 $X=284550 $Y=323440
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 345440 1 0 $X=298810 $Y=342480
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=301760 312800 0 0 $X=301570 $Y=312560
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=310960 318240 0 0 $X=310770 $Y=318000
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=313260 312800 1 0 $X=313070 $Y=309840
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=317400 329120 1 0 $X=317210 $Y=326160
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=347760 329120 1 0 $X=347570 $Y=326160
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=347760 350880 1 0 $X=347570 $Y=347920
X78 1 2 ICV_1 $T=5520 312800 1 0 $X=5330 $Y=309840
X79 1 2 ICV_1 $T=5520 318240 1 0 $X=5330 $Y=315280
X80 1 2 ICV_1 $T=5520 323680 1 0 $X=5330 $Y=320720
X81 1 2 ICV_1 $T=5520 329120 1 0 $X=5330 $Y=326160
X82 1 2 ICV_1 $T=5520 334560 1 0 $X=5330 $Y=331600
X83 1 2 ICV_1 $T=5520 340000 1 0 $X=5330 $Y=337040
X84 1 2 ICV_1 $T=5520 345440 1 0 $X=5330 $Y=342480
X85 1 2 ICV_1 $T=5520 350880 1 0 $X=5330 $Y=347920
X86 1 2 ICV_1 $T=350520 312800 0 180 $X=348950 $Y=309840
X87 1 2 ICV_1 $T=350520 318240 0 180 $X=348950 $Y=315280
X88 1 2 ICV_1 $T=350520 323680 0 180 $X=348950 $Y=320720
X89 1 2 ICV_1 $T=350520 329120 0 180 $X=348950 $Y=326160
X90 1 2 ICV_1 $T=350520 334560 0 180 $X=348950 $Y=331600
X91 1 2 ICV_1 $T=350520 340000 0 180 $X=348950 $Y=337040
X92 1 2 ICV_1 $T=350520 345440 0 180 $X=348950 $Y=342480
X93 1 2 ICV_1 $T=350520 350880 0 180 $X=348950 $Y=347920
X157 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 329120 0 0 $X=6710 $Y=328880
X158 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 323680 1 0 $X=15910 $Y=320720
X159 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 350880 1 0 $X=15910 $Y=347920
X160 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=31740 318240 1 0 $X=31550 $Y=315280
X161 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=31740 323680 1 0 $X=31550 $Y=320720
X162 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34040 329120 0 0 $X=33850 $Y=328880
X163 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=37260 329120 1 0 $X=37070 $Y=326160
X164 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=37260 334560 1 0 $X=37070 $Y=331600
X165 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=37720 340000 1 0 $X=37530 $Y=337040
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39560 323680 0 0 $X=39370 $Y=323440
X167 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=51060 340000 0 0 $X=50870 $Y=339760
X168 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=59800 350880 1 0 $X=59610 $Y=347920
X169 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=61180 334560 1 0 $X=60990 $Y=331600
X170 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=67620 340000 0 0 $X=67430 $Y=339760
X171 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=83720 329120 1 0 $X=83530 $Y=326160
X172 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=86020 329120 0 0 $X=85830 $Y=328880
X173 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 318240 1 0 $X=100090 $Y=315280
X174 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 334560 1 0 $X=100090 $Y=331600
X175 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 345440 1 0 $X=104230 $Y=342480
X176 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 350880 1 0 $X=104230 $Y=347920
X177 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=110860 318240 1 0 $X=110670 $Y=315280
X178 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=111320 312800 1 0 $X=111130 $Y=309840
X179 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=124660 312800 0 0 $X=124470 $Y=312560
X180 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126960 350880 1 0 $X=126770 $Y=347920
X181 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=127880 323680 1 0 $X=127690 $Y=320720
X182 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 312800 1 0 $X=128150 $Y=309840
X183 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=135240 340000 0 0 $X=135050 $Y=339760
X184 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=137540 334560 0 0 $X=137350 $Y=334320
X185 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=138000 345440 1 0 $X=137810 $Y=342480
X186 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=140760 318240 0 0 $X=140570 $Y=318000
X187 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 312800 1 0 $X=146090 $Y=309840
X188 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 312800 0 0 $X=146090 $Y=312560
X189 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 318240 0 0 $X=146090 $Y=318000
X190 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 340000 0 0 $X=146090 $Y=339760
X191 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=147660 318240 1 0 $X=147470 $Y=315280
X192 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 340000 1 0 $X=156210 $Y=337040
X193 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=160540 329120 1 0 $X=160350 $Y=326160
X194 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=161460 334560 0 0 $X=161270 $Y=334320
X195 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=163300 345440 0 0 $X=163110 $Y=345200
X196 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=166060 350880 1 0 $X=165870 $Y=347920
X197 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 312800 0 0 $X=170010 $Y=312560
X198 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=179860 340000 0 0 $X=179670 $Y=339760
X199 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=179860 345440 0 0 $X=179670 $Y=345200
X200 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=180780 312800 1 0 $X=180590 $Y=309840
X201 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=196880 334560 0 0 $X=196690 $Y=334320
X202 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198260 323680 0 0 $X=198070 $Y=323440
X203 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=200560 340000 1 0 $X=200370 $Y=337040
X204 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=202400 323680 0 0 $X=202210 $Y=323440
X205 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=204700 329120 1 0 $X=204510 $Y=326160
X206 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=214820 340000 0 0 $X=214630 $Y=339760
X207 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 340000 1 0 $X=216470 $Y=337040
X208 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=224480 340000 0 0 $X=224290 $Y=339760
X209 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239200 340000 1 0 $X=239010 $Y=337040
X210 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 334560 1 0 $X=240390 $Y=331600
X211 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=242880 329120 0 0 $X=242690 $Y=328880
X212 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=243340 323680 0 0 $X=243150 $Y=323440
X213 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=247480 334560 0 0 $X=247290 $Y=334320
X214 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254380 334560 0 0 $X=254190 $Y=334320
X215 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=256680 329120 1 0 $X=256490 $Y=326160
X216 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=264040 345440 0 0 $X=263850 $Y=345200
X217 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=270020 340000 0 0 $X=269830 $Y=339760
X218 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281520 329120 0 0 $X=281330 $Y=328880
X219 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281980 318240 0 0 $X=281790 $Y=318000
X220 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286580 318240 0 0 $X=286390 $Y=318000
X221 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=295320 345440 1 0 $X=295130 $Y=342480
X222 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=295780 318240 1 0 $X=295590 $Y=315280
X223 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=295780 350880 1 0 $X=295590 $Y=347920
X224 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 323680 1 0 $X=296510 $Y=320720
X225 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 329120 1 0 $X=296510 $Y=326160
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 334560 0 0 $X=310310 $Y=334320
X227 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=319700 318240 0 0 $X=319510 $Y=318000
X228 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=323840 318240 1 0 $X=323650 $Y=315280
X229 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324300 350880 1 0 $X=324110 $Y=347920
X230 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 312800 1 0 $X=324570 $Y=309840
X231 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 350880 1 0 $X=328710 $Y=347920
X232 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=330740 334560 0 0 $X=330550 $Y=334320
X233 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=338100 323680 0 0 $X=337910 $Y=323440
X234 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344080 350880 1 0 $X=343890 $Y=347920
X235 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 334560 1 0 $X=345270 $Y=331600
X236 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 340000 1 0 $X=345270 $Y=337040
X237 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 350880 0 0 $X=6710 $Y=350640
X238 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=42320 345440 1 0 $X=42130 $Y=342480
X239 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=75900 334560 0 0 $X=75710 $Y=334320
X240 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=80500 329120 0 0 $X=80310 $Y=328880
X241 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82800 323680 1 0 $X=82610 $Y=320720
X242 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=98440 323680 1 0 $X=98250 $Y=320720
X243 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=106720 323680 0 0 $X=106530 $Y=323440
X244 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 345440 1 0 $X=125390 $Y=342480
X245 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=135240 318240 0 0 $X=135050 $Y=318000
X246 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=165600 323680 1 0 $X=165410 $Y=320720
X247 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=179400 323680 1 0 $X=179210 $Y=320720
X248 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=191360 334560 0 0 $X=191170 $Y=334320
X249 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=191820 318240 0 0 $X=191630 $Y=318000
X250 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195040 318240 1 0 $X=194850 $Y=315280
X251 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=206080 334560 1 0 $X=205890 $Y=331600
X252 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=233680 340000 1 0 $X=233490 $Y=337040
X253 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237820 312800 1 0 $X=237630 $Y=309840
X254 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237820 318240 1 0 $X=237630 $Y=315280
X255 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237820 323680 0 0 $X=237630 $Y=323440
X256 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=238740 329120 1 0 $X=238550 $Y=326160
X257 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=263120 334560 1 0 $X=262930 $Y=331600
X258 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=279220 323680 0 0 $X=279030 $Y=323440
X259 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=306360 329120 1 0 $X=306170 $Y=326160
X260 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=311880 329120 1 0 $X=311690 $Y=326160
X261 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=312800 318240 1 0 $X=312610 $Y=315280
X262 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=318320 318240 1 0 $X=318130 $Y=315280
X263 1 2 ICV_2 $T=19780 340000 1 0 $X=19590 $Y=337040
X264 1 2 ICV_2 $T=33580 323680 0 0 $X=33390 $Y=323440
X265 1 2 ICV_2 $T=33580 334560 0 0 $X=33390 $Y=334320
X266 1 2 ICV_2 $T=47840 340000 1 0 $X=47650 $Y=337040
X267 1 2 ICV_2 $T=47840 345440 1 0 $X=47650 $Y=342480
X268 1 2 ICV_2 $T=61640 340000 0 0 $X=61450 $Y=339760
X269 1 2 ICV_2 $T=75900 312800 1 0 $X=75710 $Y=309840
X270 1 2 ICV_2 $T=103960 323680 1 0 $X=103770 $Y=320720
X271 1 2 ICV_2 $T=103960 329120 1 0 $X=103770 $Y=326160
X272 1 2 ICV_2 $T=117760 334560 0 0 $X=117570 $Y=334320
X273 1 2 ICV_2 $T=132020 340000 1 0 $X=131830 $Y=337040
X274 1 2 ICV_2 $T=132020 345440 1 0 $X=131830 $Y=342480
X275 1 2 ICV_2 $T=160080 340000 1 0 $X=159890 $Y=337040
X276 1 2 ICV_2 $T=160080 345440 1 0 $X=159890 $Y=342480
X277 1 2 ICV_2 $T=160080 350880 1 0 $X=159890 $Y=347920
X278 1 2 ICV_2 $T=173880 340000 0 0 $X=173690 $Y=339760
X279 1 2 ICV_2 $T=173880 345440 0 0 $X=173690 $Y=345200
X280 1 2 ICV_2 $T=188140 312800 1 0 $X=187950 $Y=309840
X281 1 2 ICV_2 $T=188140 329120 1 0 $X=187950 $Y=326160
X282 1 2 ICV_2 $T=201940 334560 0 0 $X=201750 $Y=334320
X283 1 2 ICV_2 $T=216200 345440 1 0 $X=216010 $Y=342480
X284 1 2 ICV_2 $T=216200 350880 1 0 $X=216010 $Y=347920
X285 1 2 ICV_2 $T=244260 323680 1 0 $X=244070 $Y=320720
X286 1 2 ICV_2 $T=244260 329120 1 0 $X=244070 $Y=326160
X287 1 2 ICV_2 $T=244260 340000 1 0 $X=244070 $Y=337040
X288 1 2 ICV_2 $T=258060 334560 0 0 $X=257870 $Y=334320
X289 1 2 ICV_2 $T=258060 345440 0 0 $X=257870 $Y=345200
X290 1 2 ICV_2 $T=286120 329120 0 0 $X=285930 $Y=328880
X291 1 2 ICV_2 $T=300380 323680 1 0 $X=300190 $Y=320720
X292 1 2 ICV_2 $T=300380 329120 1 0 $X=300190 $Y=326160
X293 1 2 ICV_2 $T=300380 350880 1 0 $X=300190 $Y=347920
X294 1 2 ICV_2 $T=328440 334560 1 0 $X=328250 $Y=331600
X295 1 2 ICV_2 $T=342240 312800 0 0 $X=342050 $Y=312560
X296 1 2 ICV_2 $T=342240 318240 0 0 $X=342050 $Y=318000
X297 1 2 ICV_2 $T=342240 323680 0 0 $X=342050 $Y=323440
X298 1 2 ICV_2 $T=342240 329120 0 0 $X=342050 $Y=328880
X299 1 2 ICV_2 $T=342240 334560 0 0 $X=342050 $Y=334320
X300 1 2 ICV_2 $T=342240 340000 0 0 $X=342050 $Y=339760
X301 1 2 ICV_2 $T=342240 345440 0 0 $X=342050 $Y=345200
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=10580 334560 1 0 $X=10390 $Y=331600
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 312800 1 0 $X=17750 $Y=309840
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 318240 1 0 $X=17750 $Y=315280
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 312800 0 0 $X=18210 $Y=312560
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 323680 0 0 $X=18210 $Y=323440
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 345440 0 0 $X=18210 $Y=345200
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=20700 340000 0 0 $X=20510 $Y=339760
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 350880 1 0 $X=31550 $Y=347920
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 318240 0 0 $X=45810 $Y=318000
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=53820 345440 1 0 $X=53630 $Y=342480
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=55660 323680 0 0 $X=55470 $Y=323440
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=57500 312800 0 0 $X=57310 $Y=312560
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=57500 318240 0 0 $X=57310 $Y=318000
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59800 329120 1 0 $X=59610 $Y=326160
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 312800 0 0 $X=61910 $Y=312560
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 345440 0 0 $X=61910 $Y=345200
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=63940 312800 1 0 $X=63750 $Y=309840
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73600 323680 1 0 $X=73410 $Y=320720
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 340000 1 0 $X=76170 $Y=337040
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 345440 1 0 $X=76170 $Y=342480
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=84180 312800 0 0 $X=83990 $Y=312560
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87860 350880 1 0 $X=87670 $Y=347920
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=93840 329120 0 0 $X=93650 $Y=328880
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 329120 0 0 $X=101930 $Y=328880
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=114080 318240 0 0 $X=113890 $Y=318000
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 323680 0 0 $X=115730 $Y=323440
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 334560 0 0 $X=115730 $Y=334320
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143980 350880 1 0 $X=143790 $Y=347920
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=152260 345440 1 0 $X=152070 $Y=342480
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 334560 1 0 $X=158050 $Y=331600
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=165140 340000 0 0 $X=164950 $Y=339760
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=166060 340000 1 0 $X=165870 $Y=337040
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 329120 1 0 $X=171850 $Y=326160
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=173420 318240 1 0 $X=173230 $Y=315280
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188140 323680 0 0 $X=187950 $Y=323440
X337 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188600 340000 1 0 $X=188410 $Y=337040
X338 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188600 345440 1 0 $X=188410 $Y=342480
X339 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=202400 340000 0 0 $X=202210 $Y=339760
X340 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=206080 345440 0 0 $X=205890 $Y=345200
X341 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=210680 340000 1 0 $X=210490 $Y=337040
X342 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=212060 312800 1 0 $X=211870 $Y=309840
X343 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 318240 1 0 $X=216470 $Y=315280
X344 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226320 312800 0 0 $X=226130 $Y=312560
X345 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226320 329120 0 0 $X=226130 $Y=328880
X346 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=228620 329120 1 0 $X=228430 $Y=326160
X347 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=234140 334560 1 0 $X=233950 $Y=331600
X348 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=240580 345440 1 0 $X=240390 $Y=342480
X349 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=240580 350880 1 0 $X=240390 $Y=347920
X350 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244720 350880 1 0 $X=244530 $Y=347920
X351 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=247020 318240 0 0 $X=246830 $Y=318000
X352 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=254380 323680 0 0 $X=254190 $Y=323440
X353 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=280140 340000 0 0 $X=279950 $Y=339760
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=282440 312800 1 0 $X=282250 $Y=309840
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=282440 345440 0 0 $X=282250 $Y=345200
X356 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=285200 329120 1 0 $X=285010 $Y=326160
X357 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286120 312800 1 0 $X=285930 $Y=309840
X358 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=293940 340000 0 0 $X=293750 $Y=339760
X359 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=300840 312800 1 0 $X=300650 $Y=309840
X360 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=306360 323680 1 0 $X=306170 $Y=320720
X361 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=308200 345440 1 0 $X=308010 $Y=342480
X362 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=312340 329120 0 0 $X=312150 $Y=328880
X363 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=322000 340000 0 0 $X=321810 $Y=339760
X364 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 323680 1 0 $X=325950 $Y=320720
X365 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=327980 312800 0 0 $X=327790 $Y=312560
X366 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 340000 1 0 $X=328710 $Y=337040
X367 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=329360 323680 0 0 $X=329170 $Y=323440
X368 1 2 ICV_3 $T=12420 350880 0 0 $X=12230 $Y=350640
X369 1 2 ICV_3 $T=40480 350880 1 0 $X=40290 $Y=347920
X370 1 2 ICV_3 $T=66700 345440 1 0 $X=66510 $Y=342480
X371 1 2 ICV_3 $T=96600 345440 1 0 $X=96410 $Y=342480
X372 1 2 ICV_3 $T=96600 350880 1 0 $X=96410 $Y=347920
X373 1 2 ICV_3 $T=101660 340000 0 0 $X=101470 $Y=339760
X374 1 2 ICV_3 $T=138000 340000 1 0 $X=137810 $Y=337040
X375 1 2 ICV_3 $T=152720 350880 1 0 $X=152530 $Y=347920
X376 1 2 ICV_3 $T=178480 340000 1 0 $X=178290 $Y=337040
X377 1 2 ICV_3 $T=180780 350880 1 0 $X=180590 $Y=347920
X378 1 2 ICV_3 $T=194120 312800 1 0 $X=193930 $Y=309840
X379 1 2 ICV_3 $T=220800 345440 0 0 $X=220610 $Y=345200
X380 1 2 ICV_3 $T=222180 345440 1 0 $X=221990 $Y=342480
X381 1 2 ICV_3 $T=222180 350880 1 0 $X=221990 $Y=347920
X382 1 2 ICV_3 $T=262660 345440 1 0 $X=262470 $Y=342480
X383 1 2 ICV_3 $T=263120 350880 1 0 $X=262930 $Y=347920
X384 1 2 ICV_3 $T=306820 323680 0 0 $X=306630 $Y=323440
X385 1 2 ICV_3 $T=320620 345440 1 0 $X=320430 $Y=342480
X386 1 2 ICV_3 $T=326140 345440 0 0 $X=325950 $Y=345200
X387 1 2 ICV_3 $T=341780 345440 1 0 $X=341590 $Y=342480
X388 1 45 sky130_fd_sc_hd__diode_2 $T=51520 318240 0 0 $X=51330 $Y=318000
X389 1 278 sky130_fd_sc_hd__diode_2 $T=57960 312800 1 0 $X=57770 $Y=309840
X390 1 53 sky130_fd_sc_hd__diode_2 $T=59800 340000 0 0 $X=59610 $Y=339760
X391 1 282 sky130_fd_sc_hd__diode_2 $T=60720 318240 1 0 $X=60530 $Y=315280
X392 1 300 sky130_fd_sc_hd__diode_2 $T=96140 329120 0 0 $X=95950 $Y=328880
X393 1 92 sky130_fd_sc_hd__diode_2 $T=119140 318240 0 0 $X=118950 $Y=318000
X394 1 75 sky130_fd_sc_hd__diode_2 $T=153640 323680 0 0 $X=153450 $Y=323440
X395 1 68 sky130_fd_sc_hd__diode_2 $T=155020 312800 0 0 $X=154830 $Y=312560
X396 1 330 sky130_fd_sc_hd__diode_2 $T=164220 329120 0 0 $X=164030 $Y=328880
X397 1 129 sky130_fd_sc_hd__diode_2 $T=172040 323680 1 0 $X=171850 $Y=320720
X398 1 4 sky130_fd_sc_hd__diode_2 $T=172040 345440 0 0 $X=171850 $Y=345200
X399 1 334 sky130_fd_sc_hd__diode_2 $T=175260 329120 0 0 $X=175070 $Y=328880
X400 1 4 sky130_fd_sc_hd__diode_2 $T=204700 318240 1 0 $X=204510 $Y=315280
X401 1 159 sky130_fd_sc_hd__diode_2 $T=218040 312800 1 0 $X=217850 $Y=309840
X402 1 349 sky130_fd_sc_hd__diode_2 $T=218500 340000 0 0 $X=218310 $Y=339760
X403 1 354 sky130_fd_sc_hd__diode_2 $T=218960 323680 1 0 $X=218770 $Y=320720
X404 1 162 sky130_fd_sc_hd__diode_2 $T=220340 329120 0 0 $X=220150 $Y=328880
X405 1 358 sky130_fd_sc_hd__diode_2 $T=229540 318240 1 0 $X=229350 $Y=315280
X406 1 75 sky130_fd_sc_hd__diode_2 $T=231840 312800 1 0 $X=231650 $Y=309840
X407 1 175 sky130_fd_sc_hd__diode_2 $T=245640 312800 0 0 $X=245450 $Y=312560
X408 1 176 sky130_fd_sc_hd__diode_2 $T=248400 323680 0 0 $X=248210 $Y=323440
X409 1 273 sky130_fd_sc_hd__diode_2 $T=250700 329120 1 0 $X=250510 $Y=326160
X410 1 370 sky130_fd_sc_hd__diode_2 $T=251160 312800 1 0 $X=250970 $Y=309840
X411 1 178 sky130_fd_sc_hd__diode_2 $T=253460 323680 1 0 $X=253270 $Y=320720
X412 1 128 sky130_fd_sc_hd__diode_2 $T=272320 312800 0 0 $X=272130 $Y=312560
X413 1 382 sky130_fd_sc_hd__diode_2 $T=300840 323680 0 0 $X=300650 $Y=323440
X414 1 2 271 ICV_4 $T=30820 334560 0 0 $X=30630 $Y=334320
X415 1 2 270 ICV_4 $T=39560 312800 1 0 $X=39370 $Y=309840
X416 1 2 274 ICV_4 $T=45080 323680 1 0 $X=44890 $Y=320720
X417 1 2 276 ICV_4 $T=50140 312800 0 0 $X=49950 $Y=312560
X418 1 2 50 ICV_4 $T=57040 329120 0 0 $X=56850 $Y=328880
X419 1 2 51 ICV_4 $T=58420 334560 0 0 $X=58230 $Y=334320
X420 1 2 282 ICV_4 $T=73140 329120 1 0 $X=72950 $Y=326160
X421 1 2 280 ICV_4 $T=97060 312800 0 0 $X=96870 $Y=312560
X422 1 2 4 ICV_4 $T=110860 345440 0 0 $X=110670 $Y=345200
X423 1 2 300 ICV_4 $T=113160 340000 0 0 $X=112970 $Y=339760
X424 1 2 93 ICV_4 $T=115000 312800 1 0 $X=114810 $Y=309840
X425 1 2 312 ICV_4 $T=133400 323680 1 0 $X=133210 $Y=320720
X426 1 2 4 ICV_4 $T=134320 329120 0 0 $X=134130 $Y=328880
X427 1 2 314 ICV_4 $T=137080 312800 1 0 $X=136890 $Y=309840
X428 1 2 311 ICV_4 $T=137080 329120 1 0 $X=136890 $Y=326160
X429 1 2 112 ICV_4 $T=141220 323680 0 0 $X=141030 $Y=323440
X430 1 2 318 ICV_4 $T=143520 323680 1 0 $X=143330 $Y=320720
X431 1 2 321 ICV_4 $T=149960 318240 0 0 $X=149770 $Y=318000
X432 1 2 324 ICV_4 $T=153640 323680 1 0 $X=153450 $Y=320720
X433 1 2 325 ICV_4 $T=156860 312800 1 0 $X=156670 $Y=309840
X434 1 2 111 ICV_4 $T=156860 318240 1 0 $X=156670 $Y=315280
X435 1 2 325 ICV_4 $T=156860 323680 1 0 $X=156670 $Y=320720
X436 1 2 118 ICV_4 $T=157320 329120 1 0 $X=157130 $Y=326160
X437 1 2 329 ICV_4 $T=162840 312800 1 0 $X=162650 $Y=309840
X438 1 2 4 ICV_4 $T=163300 312800 0 0 $X=163110 $Y=312560
X439 1 2 333 ICV_4 $T=169280 323680 0 0 $X=169090 $Y=323440
X440 1 2 4 ICV_4 $T=171120 329120 0 0 $X=170930 $Y=328880
X441 1 2 127 ICV_4 $T=171120 340000 0 0 $X=170930 $Y=339760
X442 1 2 132 ICV_4 $T=185380 318240 1 0 $X=185190 $Y=315280
X443 1 2 340 ICV_4 $T=185380 323680 1 0 $X=185190 $Y=320720
X444 1 2 345 ICV_4 $T=199180 329120 0 0 $X=198990 $Y=328880
X445 1 2 3 ICV_4 $T=199180 345440 0 0 $X=198990 $Y=345200
X446 1 2 347 ICV_4 $T=205160 323680 1 0 $X=204970 $Y=320720
X447 1 2 145 ICV_4 $T=209760 312800 0 0 $X=209570 $Y=312560
X448 1 2 153 ICV_4 $T=211600 318240 1 0 $X=211410 $Y=315280
X449 1 2 4 ICV_4 $T=212980 334560 1 0 $X=212790 $Y=331600
X450 1 2 155 ICV_4 $T=212980 340000 1 0 $X=212790 $Y=337040
X451 1 2 350 ICV_4 $T=213440 323680 1 0 $X=213250 $Y=320720
X452 1 2 357 ICV_4 $T=227240 323680 1 0 $X=227050 $Y=320720
X453 1 2 56 ICV_4 $T=231380 318240 0 0 $X=231190 $Y=318000
X454 1 2 371 ICV_4 $T=250240 323680 1 0 $X=250050 $Y=320720
X455 1 2 3 ICV_4 $T=255300 345440 0 0 $X=255110 $Y=345200
X456 1 2 180 ICV_4 $T=259440 312800 1 0 $X=259250 $Y=309840
X457 1 2 4 ICV_4 $T=269100 334560 1 0 $X=268910 $Y=331600
X458 1 2 189 ICV_4 $T=269100 340000 1 0 $X=268910 $Y=337040
X459 1 2 380 ICV_4 $T=281520 312800 0 0 $X=281330 $Y=312560
X460 1 2 199 ICV_4 $T=287960 312800 1 0 $X=287770 $Y=309840
X461 1 2 3 ICV_4 $T=311420 340000 0 0 $X=311230 $Y=339760
X462 1 2 199 ICV_4 $T=314640 312800 1 0 $X=314450 $Y=309840
X463 1 2 227 ICV_4 $T=317400 312800 1 0 $X=317210 $Y=309840
X464 1 2 4 ICV_4 $T=318780 329120 1 0 $X=318590 $Y=326160
X465 1 2 378 ICV_4 $T=339020 340000 0 0 $X=338830 $Y=339760
X466 1 2 3 ICV_4 $T=339480 318240 0 0 $X=339290 $Y=318000
X467 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 340000 1 0 $X=16370 $Y=337040
X468 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 345440 1 0 $X=16370 $Y=342480
X469 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=18400 318240 0 0 $X=18210 $Y=318000
X470 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30360 323680 0 0 $X=30170 $Y=323440
X471 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=31740 312800 1 0 $X=31550 $Y=309840
X472 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=41860 323680 1 0 $X=41670 $Y=320720
X473 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45540 345440 0 0 $X=45350 $Y=345200
X474 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=51980 334560 0 0 $X=51790 $Y=334320
X475 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=64860 329120 1 0 $X=64670 $Y=326160
X476 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 318240 0 0 $X=72950 $Y=318000
X477 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=109940 323680 1 0 $X=109750 $Y=320720
X478 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=109940 329120 1 0 $X=109750 $Y=326160
X479 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=114540 329120 0 0 $X=114350 $Y=328880
X480 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115920 340000 1 0 $X=115730 $Y=337040
X481 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=118220 329120 0 0 $X=118030 $Y=328880
X482 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=120980 312800 1 0 $X=120790 $Y=309840
X483 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129720 345440 0 0 $X=129530 $Y=345200
X484 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143980 334560 1 0 $X=143790 $Y=331600
X485 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=196880 340000 0 0 $X=196690 $Y=339760
X486 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=201020 345440 1 0 $X=200830 $Y=342480
X487 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=207000 350880 1 0 $X=206810 $Y=347920
X488 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=207920 334560 0 0 $X=207730 $Y=334320
X489 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=228160 334560 1 0 $X=227970 $Y=331600
X490 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 312800 1 0 $X=244530 $Y=309840
X491 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=264040 334560 0 0 $X=263850 $Y=334320
X492 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=264500 329120 1 0 $X=264310 $Y=326160
X493 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=278300 312800 0 0 $X=278110 $Y=312560
X494 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=283360 334560 0 0 $X=283170 $Y=334320
X495 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=284280 323680 1 0 $X=284090 $Y=320720
X496 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=284280 350880 1 0 $X=284090 $Y=347920
X497 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297160 340000 1 0 $X=296970 $Y=337040
X498 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=298080 323680 0 0 $X=297890 $Y=323440
X499 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=305440 318240 0 0 $X=305250 $Y=318000
X500 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=305900 318240 1 0 $X=305710 $Y=315280
X501 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=306360 329120 0 0 $X=306170 $Y=328880
X502 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=308200 334560 1 0 $X=308010 $Y=331600
X503 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=328900 329120 1 0 $X=328710 $Y=326160
X504 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=332120 329120 0 0 $X=331930 $Y=328880
X505 1 2 24 ICV_5 $T=26220 340000 0 0 $X=26030 $Y=339760
X506 1 2 4 ICV_5 $T=41860 329120 1 0 $X=41670 $Y=326160
X507 1 2 4 ICV_5 $T=90160 340000 1 0 $X=89970 $Y=337040
X508 1 2 301 ICV_5 $T=97980 312800 1 0 $X=97790 $Y=309840
X509 1 2 310 ICV_5 $T=122820 334560 1 0 $X=122630 $Y=331600
X510 1 2 309 ICV_5 $T=124660 329120 1 0 $X=124470 $Y=326160
X511 1 2 308 ICV_5 $T=128340 329120 1 0 $X=128150 $Y=326160
X512 1 2 109 ICV_5 $T=133400 312800 1 0 $X=133210 $Y=309840
X513 1 2 92 ICV_5 $T=133400 318240 1 0 $X=133210 $Y=315280
X514 1 2 313 ICV_5 $T=133400 329120 1 0 $X=133210 $Y=326160
X515 1 2 316 ICV_5 $T=136160 323680 1 0 $X=135970 $Y=320720
X516 1 2 336 ICV_5 $T=174340 329120 1 0 $X=174150 $Y=326160
X517 1 2 337 ICV_5 $T=175260 312800 0 0 $X=175070 $Y=312560
X518 1 2 339 ICV_5 $T=184000 329120 1 0 $X=183810 $Y=326160
X519 1 2 355 ICV_5 $T=225860 318240 1 0 $X=225670 $Y=315280
X520 1 2 177 ICV_5 $T=252080 340000 0 0 $X=251890 $Y=339760
X521 1 2 221 ICV_5 $T=310500 312800 0 0 $X=310310 $Y=312560
X522 1 2 232 ICV_5 $T=338560 329120 0 0 $X=338370 $Y=328880
X523 1 2 345 ICV_5 $T=338560 334560 0 0 $X=338370 $Y=334320
X524 1 2 4 ICV_6 $T=7820 329120 1 0 $X=7630 $Y=326160
X525 1 2 270 ICV_6 $T=23920 312800 0 0 $X=23730 $Y=312560
X526 1 2 22 ICV_6 $T=27600 329120 0 0 $X=27410 $Y=328880
X527 1 2 40 ICV_6 $T=42320 312800 1 0 $X=42130 $Y=309840
X528 1 2 4 ICV_6 $T=65320 334560 1 0 $X=65130 $Y=331600
X529 1 2 287 ICV_6 $T=69920 334560 1 0 $X=69730 $Y=331600
X530 1 2 290 ICV_6 $T=80040 323680 0 0 $X=79850 $Y=323440
X531 1 2 307 ICV_6 $T=126040 318240 1 0 $X=125850 $Y=315280
X532 1 2 4 ICV_6 $T=126960 334560 1 0 $X=126770 $Y=331600
X533 1 2 105 ICV_6 $T=126960 340000 1 0 $X=126770 $Y=337040
X534 1 2 315 ICV_6 $T=136160 345440 0 0 $X=135970 $Y=345200
X535 1 2 4 ICV_6 $T=140300 312800 0 0 $X=140110 $Y=312560
X536 1 2 4 ICV_6 $T=154560 345440 1 0 $X=154370 $Y=342480
X537 1 2 343 ICV_6 $T=189520 323680 1 0 $X=189330 $Y=320720
X538 1 2 340 ICV_6 $T=192740 312800 0 0 $X=192550 $Y=312560
X539 1 2 344 ICV_6 $T=194120 323680 1 0 $X=193930 $Y=320720
X540 1 2 4 ICV_6 $T=204240 345440 1 0 $X=204050 $Y=342480
X541 1 2 4 ICV_6 $T=210220 345440 1 0 $X=210030 $Y=342480
X542 1 2 349 ICV_6 $T=210220 350880 1 0 $X=210030 $Y=347920
X543 1 2 188 ICV_6 $T=267260 312800 1 0 $X=267070 $Y=309840
X544 1 2 377 ICV_6 $T=267260 329120 1 0 $X=267070 $Y=326160
X545 1 2 4 ICV_6 $T=287500 323680 1 0 $X=287310 $Y=320720
X546 1 2 4 ICV_6 $T=290720 334560 1 0 $X=290530 $Y=331600
X547 1 2 205 ICV_6 $T=295780 334560 1 0 $X=295590 $Y=331600
X548 1 2 241 ICV_6 $T=337180 345440 0 0 $X=336990 $Y=345200
X549 1 3 4 ICV_7 $T=7820 312800 1 0 $X=7630 $Y=309840
X550 1 3 4 ICV_7 $T=7820 318240 1 0 $X=7630 $Y=315280
X551 1 3 8 ICV_7 $T=7820 334560 1 0 $X=7630 $Y=331600
X552 1 3 4 ICV_7 $T=20240 312800 0 0 $X=20050 $Y=312560
X553 1 3 4 ICV_7 $T=20240 323680 0 0 $X=20050 $Y=323440
X554 1 3 4 ICV_7 $T=20240 345440 0 0 $X=20050 $Y=345200
X555 1 3 4 ICV_7 $T=21160 318240 0 0 $X=20970 $Y=318000
X556 1 3 4 ICV_7 $T=22540 340000 0 0 $X=22350 $Y=339760
X557 1 3 4 ICV_7 $T=23920 329120 0 0 $X=23730 $Y=328880
X558 1 3 4 ICV_7 $T=27140 334560 0 0 $X=26950 $Y=334320
X559 1 272 4 ICV_7 $T=29900 312800 0 0 $X=29710 $Y=312560
X560 1 4 3 ICV_7 $T=29900 340000 0 0 $X=29710 $Y=339760
X561 1 37 3 ICV_7 $T=38180 329120 0 0 $X=37990 $Y=328880
X562 1 44 4 ICV_7 $T=46460 312800 0 0 $X=46270 $Y=312560
X563 1 275 45 ICV_7 $T=47840 318240 0 0 $X=47650 $Y=318000
X564 1 3 4 ICV_7 $T=48300 345440 0 0 $X=48110 $Y=345200
X565 1 3 4 ICV_7 $T=49220 323680 1 0 $X=49030 $Y=320720
X566 1 3 4 ICV_7 $T=53360 329120 0 0 $X=53170 $Y=328880
X567 1 277 52 ICV_7 $T=54280 312800 1 0 $X=54090 $Y=309840
X568 1 3 4 ICV_7 $T=54740 334560 0 0 $X=54550 $Y=334320
X569 1 3 4 ICV_7 $T=56120 340000 0 0 $X=55930 $Y=339760
X570 1 279 280 ICV_7 $T=57960 323680 0 0 $X=57770 $Y=323440
X571 1 279 58 ICV_7 $T=58420 323680 1 0 $X=58230 $Y=320720
X572 1 282 283 ICV_7 $T=62100 329120 1 0 $X=61910 $Y=326160
X573 1 3 4 ICV_7 $T=64400 350880 1 0 $X=64210 $Y=347920
X574 1 280 284 ICV_7 $T=70380 318240 0 0 $X=70190 $Y=318000
X575 1 288 280 ICV_7 $T=70840 323680 1 0 $X=70650 $Y=320720
X576 1 68 290 ICV_7 $T=76360 318240 0 0 $X=76170 $Y=318000
X577 1 3 4 ICV_7 $T=76360 345440 0 0 $X=76170 $Y=345200
X578 1 3 4 ICV_7 $T=78660 340000 1 0 $X=78470 $Y=337040
X579 1 292 45 ICV_7 $T=86020 312800 0 0 $X=85830 $Y=312560
X580 1 293 280 ICV_7 $T=86020 323680 0 0 $X=85830 $Y=323440
X581 1 72 3 ICV_7 $T=86020 340000 0 0 $X=85830 $Y=339760
X582 1 294 295 ICV_7 $T=87860 329120 1 0 $X=87670 $Y=326160
X583 1 295 75 ICV_7 $T=89240 323680 1 0 $X=89050 $Y=320720
X584 1 282 298 ICV_7 $T=90160 318240 1 0 $X=89970 $Y=315280
X585 1 4 297 ICV_7 $T=91080 329120 0 0 $X=90890 $Y=328880
X586 1 78 299 ICV_7 $T=94300 312800 1 0 $X=94110 $Y=309840
X587 1 299 82 ICV_7 $T=99820 312800 0 0 $X=99630 $Y=312560
X588 1 3 4 ICV_7 $T=104420 329120 0 0 $X=104230 $Y=328880
X589 1 3 4 ICV_7 $T=105800 334560 0 0 $X=105610 $Y=334320
X590 1 87 3 ICV_7 $T=107180 345440 0 0 $X=106990 $Y=345200
X591 1 89 302 ICV_7 $T=108560 312800 0 0 $X=108370 $Y=312560
X592 1 3 4 ICV_7 $T=109480 340000 0 0 $X=109290 $Y=339760
X593 1 303 91 ICV_7 $T=111320 318240 0 0 $X=111130 $Y=318000
X594 1 304 92 ICV_7 $T=112240 312800 0 0 $X=112050 $Y=312560
X595 1 4 305 ICV_7 $T=113160 323680 0 0 $X=112970 $Y=323440
X596 1 4 3 ICV_7 $T=114080 345440 0 0 $X=113890 $Y=345200
X597 1 82 304 ICV_7 $T=118220 312800 1 0 $X=118030 $Y=309840
X598 1 82 307 ICV_7 $T=118680 323680 1 0 $X=118490 $Y=320720
X599 1 101 93 ICV_7 $T=122360 318240 1 0 $X=122170 $Y=315280
X600 1 93 108 ICV_7 $T=129260 312800 0 0 $X=129070 $Y=312560
X601 1 3 4 ICV_7 $T=132480 345440 0 0 $X=132290 $Y=345200
X602 1 111 317 ICV_7 $T=139840 323680 1 0 $X=139650 $Y=320720
X603 1 311 3 ICV_7 $T=139840 340000 0 0 $X=139650 $Y=339760
X604 1 315 319 ICV_7 $T=142140 329120 0 0 $X=141950 $Y=328880
X605 1 113 4 ICV_7 $T=142140 334560 0 0 $X=141950 $Y=334320
X606 1 114 3 ICV_7 $T=142140 345440 0 0 $X=141950 $Y=345200
X607 1 118 317 ICV_7 $T=146280 323680 1 0 $X=146090 $Y=320720
X608 1 3 4 ICV_7 $T=147200 334560 0 0 $X=147010 $Y=334320
X609 1 112 111 ICV_7 $T=149960 323680 1 0 $X=149770 $Y=320720
X610 1 119 3 ICV_7 $T=150880 340000 0 0 $X=150690 $Y=339760
X611 1 320 118 ICV_7 $T=151340 312800 0 0 $X=151150 $Y=312560
X612 1 323 112 ICV_7 $T=153180 318240 0 0 $X=152990 $Y=318000
X613 1 327 328 ICV_7 $T=160540 329120 0 0 $X=160350 $Y=328880
X614 1 324 111 ICV_7 $T=161920 323680 0 0 $X=161730 $Y=323440
X615 1 123 326 ICV_7 $T=164220 318240 0 0 $X=164030 $Y=318000
X616 1 112 332 ICV_7 $T=165600 323680 0 0 $X=165410 $Y=323440
X617 1 331 3 ICV_7 $T=166060 334560 0 0 $X=165870 $Y=334320
X618 1 3 4 ICV_7 $T=167440 340000 0 0 $X=167250 $Y=339760
X619 1 332 335 ICV_7 $T=168360 318240 0 0 $X=168170 $Y=318000
X620 1 327 3 ICV_7 $T=168360 345440 0 0 $X=168170 $Y=345200
X621 1 131 132 ICV_7 $T=175260 318240 1 0 $X=175070 $Y=315280
X622 1 135 136 ICV_7 $T=178020 312800 1 0 $X=177830 $Y=309840
X623 1 101 335 ICV_7 $T=178940 312800 0 0 $X=178750 $Y=312560
X624 1 338 123 ICV_7 $T=180320 323680 0 0 $X=180130 $Y=323440
X625 1 4 3 ICV_7 $T=184000 345440 0 0 $X=183810 $Y=345200
X626 1 139 129 ICV_7 $T=189060 312800 0 0 $X=188870 $Y=312560
X627 1 4 341 ICV_7 $T=189980 329120 0 0 $X=189790 $Y=328880
X628 1 342 4 ICV_7 $T=190440 323680 0 0 $X=190250 $Y=323440
X629 1 3 4 ICV_7 $T=190440 340000 1 0 $X=190250 $Y=337040
X630 1 142 139 ICV_7 $T=198260 312800 0 0 $X=198070 $Y=312560
X631 1 346 145 ICV_7 $T=198260 318240 0 0 $X=198070 $Y=318000
X632 1 4 144 ICV_7 $T=203320 345440 0 0 $X=203130 $Y=345200
X633 1 150 154 ICV_7 $T=209300 312800 1 0 $X=209110 $Y=309840
X634 1 4 353 ICV_7 $T=216660 329120 0 0 $X=216470 $Y=328880
X635 1 352 356 ICV_7 $T=218500 329120 1 0 $X=218310 $Y=326160
X636 1 357 159 ICV_7 $T=220340 323680 0 0 $X=220150 $Y=323440
X637 1 145 351 ICV_7 $T=222180 312800 1 0 $X=221990 $Y=309840
X638 1 57 165 ICV_7 $T=224020 318240 0 0 $X=223830 $Y=318000
X639 1 3 4 ICV_7 $T=224480 334560 0 0 $X=224290 $Y=334320
X640 1 358 159 ICV_7 $T=226320 323680 0 0 $X=226130 $Y=323440
X641 1 359 168 ICV_7 $T=228160 312800 1 0 $X=227970 $Y=309840
X642 1 4 362 ICV_7 $T=231380 334560 1 0 $X=231190 $Y=331600
X643 1 157 165 ICV_7 $T=238280 312800 0 0 $X=238090 $Y=312560
X644 1 4 3 ICV_7 $T=240120 345440 0 0 $X=239930 $Y=345200
X645 1 365 366 ICV_7 $T=241960 312800 0 0 $X=241770 $Y=312560
X646 1 165 370 ICV_7 $T=247480 312800 1 0 $X=247290 $Y=309840
X647 1 3 4 ICV_7 $T=248400 340000 0 0 $X=248210 $Y=339760
X648 1 369 367 ICV_7 $T=248860 318240 0 0 $X=248670 $Y=318000
X649 1 4 372 ICV_7 $T=251620 334560 0 0 $X=251430 $Y=334320
X650 1 366 180 ICV_7 $T=252540 318240 0 0 $X=252350 $Y=318000
X651 1 3 289 ICV_7 $T=259900 345440 1 0 $X=259710 $Y=342480
X652 1 178 183 ICV_7 $T=260820 318240 1 0 $X=260630 $Y=315280
X653 1 3 3 ICV_7 $T=268180 345440 0 0 $X=267990 $Y=345200
X654 1 4 4 ICV_7 $T=273700 345440 1 0 $X=273510 $Y=342480
X655 1 3 4 ICV_7 $T=278760 329120 0 0 $X=278570 $Y=328880
X656 1 3 4 ICV_7 $T=280600 334560 0 0 $X=280410 $Y=334320
X657 1 309 4 ICV_7 $T=282440 340000 0 0 $X=282250 $Y=339760
X658 1 296 4 ICV_7 $T=291180 318240 0 0 $X=290990 $Y=318000
X659 1 4 3 ICV_7 $T=296240 340000 0 0 $X=296050 $Y=339760
X660 1 384 199 ICV_7 $T=299000 312800 0 0 $X=298810 $Y=312560
X661 1 212 213 ICV_7 $T=303140 312800 0 0 $X=302950 $Y=312560
X662 1 214 3 ICV_7 $T=304520 345440 0 0 $X=304330 $Y=345200
X663 1 216 199 ICV_7 $T=306820 312800 0 0 $X=306630 $Y=312560
X664 1 4 385 ICV_7 $T=308200 318240 0 0 $X=308010 $Y=318000
X665 1 218 3 ICV_7 $T=309580 329120 0 0 $X=309390 $Y=328880
X666 1 220 224 ICV_7 $T=310500 312800 1 0 $X=310310 $Y=309840
X667 1 4 3 ICV_7 $T=310500 345440 0 0 $X=310310 $Y=345200
X668 1 386 3 ICV_7 $T=316480 334560 0 0 $X=316290 $Y=334320
X669 1 320 3 ICV_7 $T=317860 329120 0 0 $X=317670 $Y=328880
X670 1 4 3 ICV_7 $T=323840 340000 0 0 $X=323650 $Y=339760
X671 1 4 3 ICV_7 $T=324300 318240 0 0 $X=324110 $Y=318000
X672 1 365 3 ICV_7 $T=330280 312800 0 0 $X=330090 $Y=312560
X673 1 3 4 ICV_7 $T=331200 340000 1 0 $X=331010 $Y=337040
X674 1 3 4 ICV_7 $T=331660 323680 0 0 $X=331470 $Y=323440
X675 1 3 4 ICV_7 $T=333500 345440 0 0 $X=333310 $Y=345200
X676 1 3 4 ICV_7 $T=334880 329120 0 0 $X=334690 $Y=328880
X677 1 3 4 ICV_7 $T=334880 334560 0 0 $X=334690 $Y=334320
X678 1 240 350 ICV_7 $T=335340 323680 0 0 $X=335150 $Y=323440
X679 1 2 3 5 4 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 312800 0 0 $X=7630 $Y=312560
X680 1 2 3 6 4 2 13 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 318240 0 0 $X=7630 $Y=318000
X681 1 2 3 7 4 2 14 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 323680 0 0 $X=7630 $Y=323440
X682 1 2 3 8 4 2 15 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 334560 0 0 $X=7630 $Y=334320
X683 1 2 3 9 4 2 16 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 345440 0 0 $X=7630 $Y=345200
X684 1 2 3 24 4 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=22540 345440 1 0 $X=22350 $Y=342480
X685 1 2 3 271 4 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=27140 340000 1 0 $X=26950 $Y=337040
X686 1 2 3 33 4 2 42 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 345440 0 0 $X=34770 $Y=345200
X687 1 2 387 31 4 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=35420 318240 0 0 $X=35230 $Y=318000
X688 1 2 3 37 4 2 49 1 sky130_fd_sc_hd__dfrtp_4 $T=41860 329120 0 0 $X=41670 $Y=328880
X689 1 2 3 43 4 2 54 1 sky130_fd_sc_hd__dfrtp_4 $T=49220 329120 1 0 $X=49030 $Y=326160
X690 1 2 3 50 4 2 59 1 sky130_fd_sc_hd__dfrtp_4 $T=50600 334560 1 0 $X=50410 $Y=331600
X691 1 2 3 51 4 2 61 1 sky130_fd_sc_hd__dfrtp_4 $T=54740 340000 1 0 $X=54550 $Y=337040
X692 1 2 3 53 4 2 63 1 sky130_fd_sc_hd__dfrtp_4 $T=56120 345440 1 0 $X=55930 $Y=342480
X693 1 2 3 281 4 2 66 1 sky130_fd_sc_hd__dfrtp_4 $T=64400 345440 0 0 $X=64210 $Y=345200
X694 1 2 3 291 4 2 74 1 sky130_fd_sc_hd__dfrtp_4 $T=78660 345440 1 0 $X=78470 $Y=342480
X695 1 2 388 70 4 2 77 1 sky130_fd_sc_hd__dfrtp_4 $T=82800 312800 1 0 $X=82610 $Y=309840
X696 1 2 389 297 4 2 300 1 sky130_fd_sc_hd__dfrtp_4 $T=89700 334560 1 0 $X=89510 $Y=331600
X697 1 2 3 87 4 2 97 1 sky130_fd_sc_hd__dfrtp_4 $T=109020 350880 1 0 $X=108830 $Y=347920
X698 1 2 390 305 4 2 309 1 sky130_fd_sc_hd__dfrtp_4 $T=113160 329120 1 0 $X=112970 $Y=326160
X699 1 2 391 314 4 2 320 1 sky130_fd_sc_hd__dfrtp_4 $T=137080 318240 1 0 $X=136890 $Y=315280
X700 1 2 3 311 4 2 120 1 sky130_fd_sc_hd__dfrtp_4 $T=141680 345440 1 0 $X=141490 $Y=342480
X701 1 2 3 113 4 2 121 1 sky130_fd_sc_hd__dfrtp_4 $T=145820 340000 1 0 $X=145630 $Y=337040
X702 1 2 392 322 4 2 327 1 sky130_fd_sc_hd__dfrtp_4 $T=150880 334560 0 0 $X=150690 $Y=334320
X703 1 2 3 119 4 2 124 1 sky130_fd_sc_hd__dfrtp_4 $T=154560 340000 0 0 $X=154370 $Y=339760
X704 1 2 393 329 4 2 126 1 sky130_fd_sc_hd__dfrtp_4 $T=162840 318240 1 0 $X=162650 $Y=315280
X705 1 2 3 127 4 2 133 1 sky130_fd_sc_hd__dfrtp_4 $T=167440 345440 1 0 $X=167250 $Y=342480
X706 1 2 3 331 4 2 134 1 sky130_fd_sc_hd__dfrtp_4 $T=167900 340000 1 0 $X=167710 $Y=337040
X707 1 2 394 330 4 2 331 1 sky130_fd_sc_hd__dfrtp_4 $T=168820 334560 1 0 $X=168630 $Y=331600
X708 1 2 3 327 4 2 137 1 sky130_fd_sc_hd__dfrtp_4 $T=170200 350880 1 0 $X=170010 $Y=347920
X709 1 2 3 342 4 2 143 1 sky130_fd_sc_hd__dfrtp_4 $T=187680 345440 0 0 $X=187490 $Y=345200
X710 1 2 3 140 4 2 147 1 sky130_fd_sc_hd__dfrtp_4 $T=190440 345440 1 0 $X=190250 $Y=342480
X711 1 2 395 344 4 2 342 1 sky130_fd_sc_hd__dfrtp_4 $T=194120 329120 1 0 $X=193930 $Y=326160
X712 1 2 3 144 4 2 152 1 sky130_fd_sc_hd__dfrtp_4 $T=196420 350880 1 0 $X=196230 $Y=347920
X713 1 2 3 146 4 2 156 1 sky130_fd_sc_hd__dfrtp_4 $T=204240 340000 0 0 $X=204050 $Y=339760
X714 1 2 396 347 4 2 158 1 sky130_fd_sc_hd__dfrtp_4 $T=204700 318240 0 0 $X=204510 $Y=318000
X715 1 2 3 166 4 2 171 1 sky130_fd_sc_hd__dfrtp_4 $T=230000 345440 1 0 $X=229810 $Y=342480
X716 1 2 3 167 4 2 172 1 sky130_fd_sc_hd__dfrtp_4 $T=230000 350880 1 0 $X=229810 $Y=347920
X717 1 2 3 173 4 2 179 1 sky130_fd_sc_hd__dfrtp_4 $T=243800 345440 0 0 $X=243610 $Y=345200
X718 1 2 3 177 4 2 185 1 sky130_fd_sc_hd__dfrtp_4 $T=248400 345440 1 0 $X=248210 $Y=342480
X719 1 2 3 289 4 2 190 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 340000 0 0 $X=259250 $Y=339760
X720 1 2 397 377 4 2 378 1 sky130_fd_sc_hd__dfrtp_4 $T=267260 329120 0 0 $X=267070 $Y=328880
X721 1 2 3 364 4 2 194 1 sky130_fd_sc_hd__dfrtp_4 $T=271860 345440 0 0 $X=271670 $Y=345200
X722 1 2 3 191 4 2 196 1 sky130_fd_sc_hd__dfrtp_4 $T=273700 350880 1 0 $X=273510 $Y=347920
X723 1 2 3 309 4 2 204 1 sky130_fd_sc_hd__dfrtp_4 $T=284740 345440 1 0 $X=284550 $Y=342480
X724 1 2 398 200 4 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=287500 312800 0 0 $X=287310 $Y=312560
X725 1 2 399 383 4 2 382 1 sky130_fd_sc_hd__dfrtp_4 $T=294860 318240 0 0 $X=294670 $Y=318000
X726 1 2 3 205 4 2 215 1 sky130_fd_sc_hd__dfrtp_4 $T=295780 329120 0 0 $X=295590 $Y=328880
X727 1 2 3 210 4 2 219 1 sky130_fd_sc_hd__dfrtp_4 $T=299920 340000 0 0 $X=299730 $Y=339760
X728 1 2 3 214 4 2 225 1 sky130_fd_sc_hd__dfrtp_4 $T=306360 350880 1 0 $X=306170 $Y=347920
X729 1 2 400 385 4 2 386 1 sky130_fd_sc_hd__dfrtp_4 $T=308200 323680 1 0 $X=308010 $Y=320720
X730 1 2 3 222 4 2 229 1 sky130_fd_sc_hd__dfrtp_4 $T=310040 345440 1 0 $X=309850 $Y=342480
X731 1 2 3 386 4 2 237 1 sky130_fd_sc_hd__dfrtp_4 $T=320160 334560 0 0 $X=319970 $Y=334320
X732 1 2 3 320 4 2 238 1 sky130_fd_sc_hd__dfrtp_4 $T=321540 329120 0 0 $X=321350 $Y=328880
X733 1 2 3 234 4 2 242 1 sky130_fd_sc_hd__dfrtp_4 $T=327520 340000 0 0 $X=327330 $Y=339760
X734 1 2 3 236 4 2 243 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 318240 0 0 $X=327790 $Y=318000
X735 1 2 3 378 4 2 244 1 sky130_fd_sc_hd__dfrtp_4 $T=331200 345440 1 0 $X=331010 $Y=342480
X736 1 2 3 241 4 2 249 1 sky130_fd_sc_hd__dfrtp_4 $T=333500 350880 1 0 $X=333310 $Y=347920
X737 1 2 3 232 4 2 250 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 334560 1 0 $X=334690 $Y=331600
X738 1 2 3 345 4 2 251 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 340000 1 0 $X=334690 $Y=337040
X739 1 2 3 7 ICV_8 $T=7820 323680 1 0 $X=7630 $Y=320720
X740 1 2 4 9 ICV_8 $T=7820 350880 1 0 $X=7630 $Y=347920
X741 1 2 4 273 ICV_8 $T=34040 345440 1 0 $X=33850 $Y=342480
X742 1 2 285 64 ICV_8 $T=66240 312800 1 0 $X=66050 $Y=309840
X743 1 2 4 79 ICV_8 $T=94300 340000 1 0 $X=94110 $Y=337040
X744 1 2 282 76 ICV_8 $T=98440 323680 0 0 $X=98250 $Y=323440
X745 1 2 3 99 ICV_8 $T=118680 340000 1 0 $X=118490 $Y=337040
X746 1 2 125 126 ICV_8 $T=166060 312800 1 0 $X=165870 $Y=309840
X747 1 2 157 361 ICV_8 $T=230460 329120 1 0 $X=230270 $Y=326160
X748 1 2 3 4 ICV_8 $T=231380 340000 0 0 $X=231190 $Y=339760
X749 1 2 3 4 ICV_8 $T=231380 345440 0 0 $X=231190 $Y=345200
X750 1 2 4 368 ICV_8 $T=247020 329120 0 0 $X=246830 $Y=328880
X751 1 2 176 374 ICV_8 $T=262660 323680 1 0 $X=262470 $Y=320720
X752 1 2 373 375 ICV_8 $T=264500 323680 0 0 $X=264310 $Y=323440
X753 1 2 4 379 ICV_8 $T=273700 318240 0 0 $X=273510 $Y=318000
X754 1 2 3 201 ICV_8 $T=287500 350880 1 0 $X=287310 $Y=347920
X755 1 2 3 4 ICV_8 $T=302220 334560 0 0 $X=302030 $Y=334320
X756 1 2 4 239 ICV_8 $T=333960 312800 0 0 $X=333770 $Y=312560
X757 1 2 ICV_9 $T=18400 334560 0 0 $X=18210 $Y=334320
X758 1 2 ICV_9 $T=39560 318240 1 0 $X=39370 $Y=315280
X759 1 2 ICV_9 $T=67160 350880 1 0 $X=66970 $Y=347920
X760 1 2 ICV_9 $T=81420 318240 1 0 $X=81230 $Y=315280
X761 1 2 ICV_9 $T=81420 334560 1 0 $X=81230 $Y=331600
X762 1 2 ICV_9 $T=81420 334560 0 0 $X=81230 $Y=334320
X763 1 2 ICV_9 $T=95680 329120 1 0 $X=95490 $Y=326160
X764 1 2 ICV_9 $T=151800 329120 0 0 $X=151610 $Y=328880
X765 1 2 ICV_9 $T=178020 345440 1 0 $X=177830 $Y=342480
X766 1 2 ICV_9 $T=179400 334560 1 0 $X=179210 $Y=331600
X767 1 2 ICV_9 $T=239660 340000 0 0 $X=239470 $Y=339760
X768 1 2 ICV_9 $T=276460 345440 1 0 $X=276270 $Y=342480
X769 1 2 ICV_10 $T=201940 329120 0 0 $X=201750 $Y=328880
X770 1 2 ICV_10 $T=333500 350880 0 0 $X=333310 $Y=350640
X771 1 2 3 20 28 4 ICV_11 $T=21160 329120 1 0 $X=20970 $Y=326160
X772 1 2 3 22 29 4 ICV_11 $T=21160 334560 1 0 $X=20970 $Y=331600
X773 1 2 3 273 41 4 ICV_11 $T=34960 340000 0 0 $X=34770 $Y=339760
X774 1 2 3 296 81 4 ICV_11 $T=91080 345440 0 0 $X=90890 $Y=345200
X775 1 2 401 298 83 4 ICV_11 $T=93840 318240 0 0 $X=93650 $Y=318000
X776 1 2 3 77 94 4 ICV_11 $T=105340 334560 1 0 $X=105150 $Y=331600
X777 1 2 3 300 98 4 ICV_11 $T=109480 345440 1 0 $X=109290 $Y=342480
X778 1 2 3 99 106 4 ICV_11 $T=119140 340000 0 0 $X=118950 $Y=339760
X779 1 2 3 114 122 4 ICV_11 $T=147200 345440 0 0 $X=147010 $Y=345200
X780 1 2 402 334 338 4 ICV_11 $T=175260 334560 0 0 $X=175070 $Y=334320
X781 1 2 403 341 345 4 ICV_11 $T=189980 334560 1 0 $X=189790 $Y=331600
X782 1 2 404 360 364 4 ICV_11 $T=231380 334560 0 0 $X=231190 $Y=334320
X783 1 2 405 368 273 4 ICV_11 $T=247020 334560 1 0 $X=246830 $Y=331600
X784 1 2 3 174 184 4 ICV_11 $T=247020 350880 1 0 $X=246830 $Y=347920
X785 1 2 406 372 281 4 ICV_11 $T=251620 340000 1 0 $X=251430 $Y=337040
X786 1 2 3 338 195 4 ICV_11 $T=273700 340000 1 0 $X=273510 $Y=337040
X787 1 2 3 380 197 4 ICV_11 $T=274620 334560 1 0 $X=274430 $Y=331600
X788 1 2 3 201 207 4 ICV_11 $T=287500 345440 0 0 $X=287310 $Y=345200
X789 1 2 3 218 231 4 ICV_11 $T=311420 334560 1 0 $X=311230 $Y=331600
X790 1 2 3 350 245 4 ICV_11 $T=331660 329120 1 0 $X=331470 $Y=326160
X791 1 2 3 365 246 4 ICV_11 $T=332120 318240 1 0 $X=331930 $Y=315280
X792 1 2 3 239 247 4 ICV_11 $T=332580 312800 1 0 $X=332390 $Y=309840
X793 1 2 3 240 248 4 ICV_11 $T=332580 323680 1 0 $X=332390 $Y=320720
X794 1 2 4 ICV_12 $T=7820 340000 1 0 $X=7630 $Y=337040
X795 1 2 3 ICV_12 $T=7820 345440 1 0 $X=7630 $Y=342480
X796 1 2 286 ICV_12 $T=68540 323680 1 0 $X=68350 $Y=320720
X797 1 2 45 ICV_12 $T=70380 323680 0 0 $X=70190 $Y=323440
X798 1 2 88 ICV_12 $T=107640 312800 1 0 $X=107450 $Y=309840
X799 1 2 4 ICV_12 $T=143520 340000 0 0 $X=143330 $Y=339760
X800 1 2 102 ICV_12 $T=147660 329120 1 0 $X=147470 $Y=326160
X801 1 2 123 ICV_12 $T=166520 334560 1 0 $X=166330 $Y=331600
X802 1 2 4 ICV_12 $T=169740 334560 0 0 $X=169550 $Y=334320
X803 1 2 135 ICV_12 $T=185840 312800 1 0 $X=185650 $Y=309840
X804 1 2 157 ICV_12 $T=224020 323680 0 0 $X=223830 $Y=323440
X805 1 2 165 ICV_12 $T=225860 312800 1 0 $X=225670 $Y=309840
X806 1 2 180 ICV_12 $T=253920 312800 0 0 $X=253730 $Y=312560
X807 1 2 5 ICV_12 $T=296240 312800 1 0 $X=296050 $Y=309840
X808 1 2 4 ICV_12 $T=308200 345440 0 0 $X=308010 $Y=345200
X809 1 2 4 ICV_12 $T=315560 329120 0 0 $X=315370 $Y=328880
X810 1 2 236 ICV_12 $T=329820 318240 1 0 $X=329630 $Y=315280
X811 1 2 4 ICV_13 $T=90160 318240 0 0 $X=89970 $Y=318000
X812 1 2 91 ICV_13 $T=124660 323680 0 0 $X=124470 $Y=323440
X813 1 2 91 ICV_13 $T=127420 318240 0 0 $X=127230 $Y=318000
X814 1 2 102 ICV_13 $T=132480 323680 0 0 $X=132290 $Y=323440
X815 1 2 131 ICV_13 $T=181700 318240 0 0 $X=181510 $Y=318000
X816 1 2 148 ICV_13 $T=200560 318240 1 0 $X=200370 $Y=315280
X817 1 2 145 ICV_13 $T=215280 318240 0 0 $X=215090 $Y=318000
X818 1 2 68 ICV_13 $T=217120 312800 0 0 $X=216930 $Y=312560
X819 1 2 4 ICV_13 $T=244720 345440 1 0 $X=244530 $Y=342480
X820 1 2 178 ICV_13 $T=249780 318240 1 0 $X=249590 $Y=315280
X821 1 2 4 ICV_13 $T=263580 329120 0 0 $X=263390 $Y=328880
X822 1 2 3 ICV_13 $T=292100 329120 0 0 $X=291910 $Y=328880
X823 1 2 383 ICV_13 $T=293020 318240 1 0 $X=292830 $Y=315280
X824 1 2 4 ICV_13 $T=293940 329120 1 0 $X=293750 $Y=326160
X825 1 2 4 ICV_13 $T=328900 312800 1 0 $X=328710 $Y=309840
X826 1 2 4 ICV_13 $T=328900 323680 1 0 $X=328710 $Y=320720
X827 1 2 ICV_14 $T=19780 345440 1 0 $X=19590 $Y=342480
X828 1 2 ICV_14 $T=47840 334560 1 0 $X=47650 $Y=331600
X829 1 2 ICV_14 $T=89700 312800 0 0 $X=89510 $Y=312560
X830 1 2 ICV_14 $T=89700 334560 0 0 $X=89510 $Y=334320
X831 1 2 ICV_14 $T=117760 323680 0 0 $X=117570 $Y=323440
X832 1 2 ICV_14 $T=160080 312800 1 0 $X=159890 $Y=309840
X833 1 2 ICV_14 $T=160080 318240 1 0 $X=159890 $Y=315280
X834 1 2 ICV_14 $T=201940 318240 0 0 $X=201750 $Y=318000
X835 1 2 ICV_14 $T=216200 323680 1 0 $X=216010 $Y=320720
X836 1 2 ICV_14 $T=216200 329120 1 0 $X=216010 $Y=326160
X837 1 2 ICV_14 $T=244260 334560 1 0 $X=244070 $Y=331600
X838 1 2 ICV_14 $T=272320 334560 1 0 $X=272130 $Y=331600
X839 1 2 ICV_14 $T=286120 334560 0 0 $X=285930 $Y=334320
X840 1 2 ICV_14 $T=314180 323680 0 0 $X=313990 $Y=323440
X841 1 2 ICV_14 $T=314180 334560 0 0 $X=313990 $Y=334320
X842 1 2 ICV_14 $T=328440 345440 1 0 $X=328250 $Y=342480
X843 1 31 ICV_15 $T=31740 318240 0 0 $X=31550 $Y=318000
X844 1 3 ICV_15 $T=31740 345440 0 0 $X=31550 $Y=345200
X845 1 43 ICV_15 $T=46000 329120 1 0 $X=45810 $Y=326160
X846 1 57 ICV_15 $T=59800 312800 0 0 $X=59610 $Y=312560
X847 1 56 ICV_15 $T=59800 318240 0 0 $X=59610 $Y=318000
X848 1 271 ICV_15 $T=59800 329120 0 0 $X=59610 $Y=328880
X849 1 281 ICV_15 $T=59800 345440 0 0 $X=59610 $Y=345200
X850 1 4 ICV_15 $T=74060 340000 1 0 $X=73870 $Y=337040
X851 1 65 ICV_15 $T=74060 345440 1 0 $X=73870 $Y=342480
X852 1 58 ICV_15 $T=87860 318240 0 0 $X=87670 $Y=318000
X853 1 3 ICV_15 $T=87860 345440 0 0 $X=87670 $Y=345200
X854 1 83 ICV_15 $T=102120 312800 1 0 $X=101930 $Y=309840
X855 1 96 ICV_15 $T=115920 312800 0 0 $X=115730 $Y=312560
X856 1 306 ICV_15 $T=115920 318240 0 0 $X=115730 $Y=318000
X857 1 4 ICV_15 $T=115920 340000 0 0 $X=115730 $Y=339760
X858 1 56 ICV_15 $T=143980 323680 0 0 $X=143790 $Y=323440
X859 1 89 ICV_15 $T=172040 318240 0 0 $X=171850 $Y=318000
X860 1 128 ICV_15 $T=172040 323680 0 0 $X=171850 $Y=323440
X861 1 4 ICV_15 $T=172040 334560 0 0 $X=171850 $Y=334320
X862 1 4 ICV_15 $T=186300 340000 1 0 $X=186110 $Y=337040
X863 1 138 ICV_15 $T=186300 345440 1 0 $X=186110 $Y=342480
X864 1 146 ICV_15 $T=200100 340000 0 0 $X=199910 $Y=339760
X865 1 157 ICV_15 $T=214360 312800 1 0 $X=214170 $Y=309840
X866 1 351 ICV_15 $T=214360 318240 1 0 $X=214170 $Y=315280
X867 1 159 ICV_15 $T=228160 312800 0 0 $X=227970 $Y=312560
X868 1 165 ICV_15 $T=228160 318240 0 0 $X=227970 $Y=318000
X869 1 145 ICV_15 $T=228160 329120 0 0 $X=227970 $Y=328880
X870 1 360 ICV_15 $T=228160 334560 0 0 $X=227970 $Y=334320
X871 1 166 ICV_15 $T=228160 340000 0 0 $X=227970 $Y=339760
X872 1 167 ICV_15 $T=228160 345440 0 0 $X=227970 $Y=345200
X873 1 174 ICV_15 $T=242420 345440 1 0 $X=242230 $Y=342480
X874 1 173 ICV_15 $T=242420 350880 1 0 $X=242230 $Y=347920
X875 1 182 ICV_15 $T=256220 312800 0 0 $X=256030 $Y=312560
X876 1 180 ICV_15 $T=256220 318240 0 0 $X=256030 $Y=318000
X877 1 162 ICV_15 $T=256220 323680 0 0 $X=256030 $Y=323440
X878 1 281 ICV_15 $T=256220 329120 0 0 $X=256030 $Y=328880
X879 1 4 ICV_15 $T=256220 340000 0 0 $X=256030 $Y=339760
X880 1 364 ICV_15 $T=270480 345440 1 0 $X=270290 $Y=342480
X881 1 191 ICV_15 $T=270480 350880 1 0 $X=270290 $Y=347920
X882 1 4 ICV_15 $T=284280 312800 0 0 $X=284090 $Y=312560
X883 1 4 ICV_15 $T=284280 345440 0 0 $X=284090 $Y=345200
X884 1 208 ICV_15 $T=298540 312800 1 0 $X=298350 $Y=309840
X885 1 386 ICV_15 $T=312340 318240 0 0 $X=312150 $Y=318000
X886 1 234 ICV_15 $T=326600 340000 1 0 $X=326410 $Y=337040
X887 1 2 4 ICV_16 $T=10120 340000 1 0 $X=9930 $Y=337040
X888 1 2 10 ICV_16 $T=10120 345440 1 0 $X=9930 $Y=342480
X889 1 2 5 ICV_16 $T=11500 312800 1 0 $X=11310 $Y=309840
X890 1 2 6 ICV_16 $T=11500 318240 1 0 $X=11310 $Y=315280
X891 1 2 4 ICV_16 $T=12420 329120 1 0 $X=12230 $Y=326160
X892 1 2 11 ICV_16 $T=12420 334560 1 0 $X=12230 $Y=331600
X893 1 2 20 ICV_16 $T=23920 323680 0 0 $X=23730 $Y=323440
X894 1 2 23 ICV_16 $T=23920 345440 0 0 $X=23730 $Y=345200
X895 1 2 19 ICV_16 $T=24840 318240 0 0 $X=24650 $Y=318000
X896 1 2 33 ICV_16 $T=34040 350880 1 0 $X=33850 $Y=347920
X897 1 2 4 ICV_16 $T=35420 323680 1 0 $X=35230 $Y=320720
X898 1 2 4 ICV_16 $T=41400 334560 1 0 $X=41210 $Y=331600
X899 1 2 39 ICV_16 $T=41400 340000 1 0 $X=41210 $Y=337040
X900 1 2 46 ICV_16 $T=51980 345440 0 0 $X=51790 $Y=345200
X901 1 2 62 ICV_16 $T=66240 340000 1 0 $X=66050 $Y=337040
X902 1 2 278 ICV_16 $T=69000 318240 1 0 $X=68810 $Y=315280
X903 1 2 291 ICV_16 $T=77280 329120 1 0 $X=77090 $Y=326160
X904 1 2 289 ICV_16 $T=77740 312800 0 0 $X=77550 $Y=312560
X905 1 2 58 ICV_16 $T=80040 318240 0 0 $X=79850 $Y=318000
X906 1 2 69 ICV_16 $T=80040 345440 0 0 $X=79850 $Y=345200
X907 1 2 291 ICV_16 $T=82340 340000 1 0 $X=82150 $Y=337040
X908 1 2 4 ICV_16 $T=90160 345440 1 0 $X=89970 $Y=342480
X909 1 2 296 ICV_16 $T=90160 350880 1 0 $X=89970 $Y=347920
X910 1 2 77 ICV_16 $T=108100 329120 0 0 $X=107910 $Y=328880
X911 1 2 86 ICV_16 $T=109480 334560 0 0 $X=109290 $Y=334320
X912 1 2 100 ICV_16 $T=120520 350880 1 0 $X=120330 $Y=347920
X913 1 2 4 ICV_16 $T=146280 350880 1 0 $X=146090 $Y=347920
X914 1 2 322 ICV_16 $T=151800 334560 1 0 $X=151610 $Y=331600
X915 1 2 331 ICV_16 $T=182160 329120 0 0 $X=181970 $Y=328880
X916 1 2 129 ICV_16 $T=182620 312800 0 0 $X=182430 $Y=312560
X917 1 2 342 ICV_16 $T=189520 350880 1 0 $X=189330 $Y=347920
X918 1 2 140 ICV_16 $T=194120 340000 1 0 $X=193930 $Y=337040
X919 1 2 3 ICV_16 $T=204240 340000 1 0 $X=204050 $Y=337040
X920 1 2 348 ICV_16 $T=208840 329120 1 0 $X=208650 $Y=326160
X921 1 2 363 ICV_16 $T=236440 323680 1 0 $X=236250 $Y=320720
X922 1 2 364 ICV_16 $T=236440 329120 0 0 $X=236250 $Y=328880
X923 1 2 376 ICV_16 $T=264500 318240 1 0 $X=264310 $Y=315280
X924 1 2 186 ICV_16 $T=265880 312800 0 0 $X=265690 $Y=312560
X925 1 2 376 ICV_16 $T=266800 318240 0 0 $X=266610 $Y=318000
X926 1 2 378 ICV_16 $T=272780 323680 0 0 $X=272590 $Y=323440
X927 1 2 338 ICV_16 $T=273700 340000 0 0 $X=273510 $Y=339760
X928 1 2 192 ICV_16 $T=274160 318240 1 0 $X=273970 $Y=315280
X929 1 2 160 ICV_16 $T=276000 312800 1 0 $X=275810 $Y=309840
X930 1 2 380 ICV_16 $T=278760 329120 1 0 $X=278570 $Y=326160
X931 1 2 200 ICV_16 $T=286580 318240 1 0 $X=286390 $Y=315280
X932 1 2 381 ICV_16 $T=287500 329120 1 0 $X=287310 $Y=326160
X933 1 2 3 ICV_16 $T=287500 340000 0 0 $X=287310 $Y=339760
X934 1 2 382 ICV_16 $T=290720 340000 1 0 $X=290530 $Y=337040
X935 1 2 211 ICV_16 $T=301760 334560 1 0 $X=301570 $Y=331600
X936 1 2 210 ICV_16 $T=301760 345440 1 0 $X=301570 $Y=342480
X937 1 2 222 ICV_16 $T=313260 340000 1 0 $X=313070 $Y=337040
X938 1 2 4 ICV_16 $T=315560 340000 0 0 $X=315370 $Y=339760
X939 1 2 226 ICV_16 $T=317860 350880 1 0 $X=317670 $Y=347920
X940 1 2 228 ICV_16 $T=319700 323680 1 0 $X=319510 $Y=320720
X941 1 2 4 ICV_16 $T=320160 340000 1 0 $X=319970 $Y=337040
X942 1 2 4 ICV_16 $T=321540 329120 1 0 $X=321350 $Y=326160
X943 1 2 270 2 38 1 sky130_fd_sc_hd__inv_8 $T=35420 318240 1 0 $X=35230 $Y=315280
X944 1 2 37 2 47 1 sky130_fd_sc_hd__inv_8 $T=49220 312800 1 0 $X=49030 $Y=309840
X945 1 2 44 2 278 1 sky130_fd_sc_hd__inv_8 $T=53360 312800 0 0 $X=53170 $Y=312560
X946 1 2 271 2 279 1 sky130_fd_sc_hd__inv_8 $T=63020 329120 0 0 $X=62830 $Y=328880
X947 1 2 289 2 64 1 sky130_fd_sc_hd__inv_8 $T=77280 318240 1 0 $X=77090 $Y=315280
X948 1 2 291 2 290 1 sky130_fd_sc_hd__inv_8 $T=77280 334560 1 0 $X=77090 $Y=331600
X949 1 2 300 2 295 1 sky130_fd_sc_hd__inv_8 $T=97980 329120 0 0 $X=97790 $Y=328880
X950 1 2 83 2 299 1 sky130_fd_sc_hd__inv_8 $T=103500 312800 0 0 $X=103310 $Y=312560
X951 1 2 309 2 304 1 sky130_fd_sc_hd__inv_8 $T=120520 323680 0 0 $X=120330 $Y=323440
X952 1 2 311 2 307 1 sky130_fd_sc_hd__inv_8 $T=137080 329120 0 0 $X=136890 $Y=328880
X953 1 2 315 2 317 1 sky130_fd_sc_hd__inv_8 $T=146740 334560 1 0 $X=146550 $Y=331600
X954 1 2 320 2 108 1 sky130_fd_sc_hd__inv_8 $T=151340 318240 1 0 $X=151150 $Y=315280
X955 1 2 327 2 324 1 sky130_fd_sc_hd__inv_8 $T=161460 334560 1 0 $X=161270 $Y=331600
X956 1 2 126 2 325 1 sky130_fd_sc_hd__inv_8 $T=166060 312800 0 0 $X=165870 $Y=312560
X957 1 2 331 2 335 1 sky130_fd_sc_hd__inv_8 $T=177100 329120 0 0 $X=176910 $Y=328880
X958 1 2 338 2 332 1 sky130_fd_sc_hd__inv_8 $T=178480 329120 1 0 $X=178290 $Y=326160
X959 1 2 342 2 142 1 sky130_fd_sc_hd__inv_8 $T=194120 323680 0 0 $X=193930 $Y=323440
X960 1 2 345 2 340 1 sky130_fd_sc_hd__inv_8 $T=194120 329120 0 0 $X=193930 $Y=328880
X961 1 2 350 2 154 1 sky130_fd_sc_hd__inv_8 $T=208380 323680 1 0 $X=208190 $Y=320720
X962 1 2 158 2 351 1 sky130_fd_sc_hd__inv_8 $T=212980 312800 0 0 $X=212790 $Y=312560
X963 1 2 349 2 357 1 sky130_fd_sc_hd__inv_8 $T=220340 340000 0 0 $X=220150 $Y=339760
X964 1 2 364 2 358 1 sky130_fd_sc_hd__inv_8 $T=236440 334560 1 0 $X=236250 $Y=331600
X965 1 2 365 2 168 1 sky130_fd_sc_hd__inv_8 $T=245640 318240 1 0 $X=245450 $Y=315280
X966 1 2 273 2 370 1 sky130_fd_sc_hd__inv_8 $T=252540 329120 1 0 $X=252350 $Y=326160
X967 1 2 281 2 376 1 sky130_fd_sc_hd__inv_8 $T=259440 329120 0 0 $X=259250 $Y=328880
X968 1 2 378 2 366 1 sky130_fd_sc_hd__inv_8 $T=273700 329120 1 0 $X=273510 $Y=326160
X969 1 2 380 2 198 1 sky130_fd_sc_hd__inv_8 $T=281520 318240 1 0 $X=281330 $Y=315280
X970 1 2 296 2 206 1 sky130_fd_sc_hd__inv_8 $T=292560 323680 1 0 $X=292370 $Y=320720
X971 1 2 382 2 213 1 sky130_fd_sc_hd__inv_8 $T=302680 323680 0 0 $X=302490 $Y=323440
X972 1 2 386 2 220 1 sky130_fd_sc_hd__inv_8 $T=315560 318240 0 0 $X=315370 $Y=318000
X973 1 2 232 2 230 1 sky130_fd_sc_hd__inv_8 $T=320620 312800 1 0 $X=320430 $Y=309840
X974 1 2 3 3 10 17 4 ICV_17 $T=8280 340000 0 0 $X=8090 $Y=339760
X975 1 2 3 3 11 21 4 ICV_17 $T=10580 329120 0 0 $X=10390 $Y=328880
X976 1 2 3 3 39 48 4 ICV_17 $T=39560 334560 0 0 $X=39370 $Y=334320
X977 1 2 4 407 274 271 4 ICV_17 $T=43240 323680 0 0 $X=43050 $Y=323440
X978 1 2 3 3 62 67 4 ICV_17 $T=63480 334560 0 0 $X=63290 $Y=334320
X979 1 2 4 408 285 289 4 ICV_17 $T=64400 312800 0 0 $X=64210 $Y=312560
X980 1 2 4 409 287 291 4 ICV_17 $T=68080 329120 0 0 $X=67890 $Y=328880
X981 1 2 3 3 65 71 4 ICV_17 $T=72220 340000 0 0 $X=72030 $Y=339760
X982 1 2 3 3 79 84 4 ICV_17 $T=92460 334560 0 0 $X=92270 $Y=334320
X983 1 2 4 410 310 311 4 ICV_17 $T=120980 329120 0 0 $X=120790 $Y=328880
X984 1 2 3 3 105 110 4 ICV_17 $T=125120 334560 0 0 $X=124930 $Y=334320
X985 1 2 3 3 138 141 4 ICV_17 $T=184460 340000 0 0 $X=184270 $Y=339760
X986 1 2 4 411 348 350 4 ICV_17 $T=207000 323680 0 0 $X=206810 $Y=323440
X987 1 2 3 3 349 161 4 ICV_17 $T=208380 345440 0 0 $X=208190 $Y=345200
X988 1 2 3 3 155 164 4 ICV_17 $T=211140 334560 0 0 $X=210950 $Y=334320
X989 1 2 163 3 163 170 4 ICV_17 $T=221260 340000 1 0 $X=221070 $Y=337040
X990 1 2 4 412 363 365 4 ICV_17 $T=234600 318240 0 0 $X=234410 $Y=318000
X991 1 2 3 3 189 193 4 ICV_17 $T=267260 334560 0 0 $X=267070 $Y=334320
X992 1 2 3 3 382 209 4 ICV_17 $T=288880 334560 0 0 $X=288690 $Y=334320
X993 1 2 4 413 227 232 4 ICV_17 $T=315560 312800 0 0 $X=315370 $Y=312560
X994 1 2 3 3 228 235 4 ICV_17 $T=316940 323680 0 0 $X=316750 $Y=323440
X995 1 2 3 18 25 4 ICV_18 $T=19780 312800 1 0 $X=19590 $Y=309840
X996 1 2 3 270 26 4 ICV_18 $T=19780 318240 1 0 $X=19590 $Y=315280
X997 1 2 3 19 27 4 ICV_18 $T=19780 323680 1 0 $X=19590 $Y=320720
X998 1 2 3 23 30 4 ICV_18 $T=19780 350880 1 0 $X=19590 $Y=347920
X999 1 2 414 272 270 4 ICV_18 $T=33580 312800 0 0 $X=33390 $Y=312560
X1000 1 2 415 276 44 4 ICV_18 $T=47840 318240 1 0 $X=47650 $Y=315280
X1001 1 2 3 46 55 4 ICV_18 $T=47840 350880 1 0 $X=47650 $Y=347920
X1002 1 2 3 69 73 4 ICV_18 $T=75900 350880 1 0 $X=75710 $Y=347920
X1003 1 2 3 72 80 4 ICV_18 $T=89700 340000 0 0 $X=89510 $Y=339760
X1004 1 2 3 86 95 4 ICV_18 $T=103960 340000 1 0 $X=103770 $Y=337040
X1005 1 2 3 100 107 4 ICV_18 $T=117760 345440 0 0 $X=117570 $Y=345200
X1006 1 2 416 313 315 4 ICV_18 $T=132020 334560 1 0 $X=131830 $Y=331600
X1007 1 2 3 315 116 4 ICV_18 $T=132020 350880 1 0 $X=131830 $Y=347920
X1008 1 2 417 353 349 4 ICV_18 $T=216200 334560 1 0 $X=216010 $Y=331600
X1009 1 2 418 379 380 4 ICV_18 $T=272320 323680 1 0 $X=272130 $Y=320720
X1010 1 2 419 381 296 4 ICV_18 $T=286120 323680 0 0 $X=285930 $Y=323440
X1011 1 2 3 211 223 4 ICV_18 $T=300380 340000 1 0 $X=300190 $Y=337040
X1012 1 2 3 226 233 4 ICV_18 $T=314180 345440 0 0 $X=313990 $Y=345200
X1013 1 2 34 35 2 272 1 sky130_fd_sc_hd__nor2_4 $T=34500 312800 1 0 $X=34310 $Y=309840
X1014 1 2 45 277 2 276 1 sky130_fd_sc_hd__nor2_4 $T=53360 318240 0 0 $X=53170 $Y=318000
X1015 1 2 45 275 2 274 1 sky130_fd_sc_hd__nor2_4 $T=53360 323680 1 0 $X=53170 $Y=320720
X1016 1 2 34 60 2 285 1 sky130_fd_sc_hd__nor2_4 $T=59800 312800 1 0 $X=59610 $Y=309840
X1017 1 2 45 286 2 287 1 sky130_fd_sc_hd__nor2_4 $T=68080 329120 1 0 $X=67890 $Y=326160
X1018 1 2 76 294 2 297 1 sky130_fd_sc_hd__nor2_4 $T=91540 329120 1 0 $X=91350 $Y=326160
X1019 1 2 45 292 2 298 1 sky130_fd_sc_hd__nor2_4 $T=92000 312800 0 0 $X=91810 $Y=312560
X1020 1 2 91 303 2 305 1 sky130_fd_sc_hd__nor2_4 $T=113160 323680 1 0 $X=112970 $Y=320720
X1021 1 2 102 103 2 104 1 sky130_fd_sc_hd__nor2_4 $T=124200 312800 1 0 $X=124010 $Y=309840
X1022 1 2 91 308 2 310 1 sky130_fd_sc_hd__nor2_4 $T=128340 323680 0 0 $X=128150 $Y=323440
X1023 1 2 91 312 2 314 1 sky130_fd_sc_hd__nor2_4 $T=131100 318240 0 0 $X=130910 $Y=318000
X1024 1 2 102 316 2 313 1 sky130_fd_sc_hd__nor2_4 $T=136160 323680 0 0 $X=135970 $Y=323440
X1025 1 2 102 319 2 322 1 sky130_fd_sc_hd__nor2_4 $T=147660 329120 0 0 $X=147470 $Y=328880
X1026 1 2 123 326 2 329 1 sky130_fd_sc_hd__nor2_4 $T=161460 323680 1 0 $X=161270 $Y=320720
X1027 1 2 123 328 2 334 1 sky130_fd_sc_hd__nor2_4 $T=166060 329120 0 0 $X=165870 $Y=328880
X1028 1 2 128 336 2 330 1 sky130_fd_sc_hd__nor2_4 $T=175260 323680 0 0 $X=175070 $Y=323440
X1029 1 2 123 339 2 341 1 sky130_fd_sc_hd__nor2_4 $T=184000 323680 0 0 $X=183810 $Y=323440
X1030 1 2 145 346 2 344 1 sky130_fd_sc_hd__nor2_4 $T=200100 323680 1 0 $X=199910 $Y=320720
X1031 1 2 145 153 2 348 1 sky130_fd_sc_hd__nor2_4 $T=206540 318240 1 0 $X=206350 $Y=315280
X1032 1 2 145 354 2 347 1 sky130_fd_sc_hd__nor2_4 $T=218960 318240 0 0 $X=218770 $Y=318000
X1033 1 2 162 352 2 353 1 sky130_fd_sc_hd__nor2_4 $T=222180 329120 0 0 $X=221990 $Y=328880
X1034 1 2 145 362 2 360 1 sky130_fd_sc_hd__nor2_4 $T=231380 329120 0 0 $X=231190 $Y=328880
X1035 1 2 162 169 2 363 1 sky130_fd_sc_hd__nor2_4 $T=233680 312800 1 0 $X=233490 $Y=309840
X1036 1 2 176 371 2 368 1 sky130_fd_sc_hd__nor2_4 $T=250240 323680 0 0 $X=250050 $Y=323440
X1037 1 2 162 373 2 377 1 sky130_fd_sc_hd__nor2_4 $T=259440 323680 0 0 $X=259250 $Y=323440
X1038 1 2 176 375 2 372 1 sky130_fd_sc_hd__nor2_4 $T=260360 329120 1 0 $X=260170 $Y=326160
X1039 1 2 162 186 2 187 1 sky130_fd_sc_hd__nor2_4 $T=262200 312800 1 0 $X=262010 $Y=309840
X1040 1 2 128 192 2 379 1 sky130_fd_sc_hd__nor2_4 $T=274160 312800 0 0 $X=273970 $Y=312560
X1041 1 2 202 203 2 381 1 sky130_fd_sc_hd__nor2_4 $T=291180 312800 1 0 $X=290990 $Y=309840
X1042 1 2 199 384 2 383 1 sky130_fd_sc_hd__nor2_4 $T=301760 318240 1 0 $X=301570 $Y=315280
X1043 1 2 199 221 2 385 1 sky130_fd_sc_hd__nor2_4 $T=308660 318240 1 0 $X=308470 $Y=315280
X1044 1 2 ICV_19 $T=19780 350880 0 0 $X=19590 $Y=350640
X1045 1 2 ICV_19 $T=48300 350880 0 0 $X=48110 $Y=350640
X1046 1 2 ICV_19 $T=76820 350880 0 0 $X=76630 $Y=350640
X1047 1 2 ICV_19 $T=105340 350880 0 0 $X=105150 $Y=350640
X1048 1 2 ICV_19 $T=133860 350880 0 0 $X=133670 $Y=350640
X1049 1 2 ICV_19 $T=162380 350880 0 0 $X=162190 $Y=350640
X1050 1 2 ICV_19 $T=190900 350880 0 0 $X=190710 $Y=350640
X1051 1 2 ICV_19 $T=219420 350880 0 0 $X=219230 $Y=350640
X1052 1 2 ICV_19 $T=247940 350880 0 0 $X=247750 $Y=350640
X1053 1 2 ICV_19 $T=276460 350880 0 0 $X=276270 $Y=350640
X1054 1 2 ICV_19 $T=304980 350880 0 0 $X=304790 $Y=350640
X1055 1 2 278 282 280 284 2 277 1 sky130_fd_sc_hd__o22a_4 $T=63020 318240 0 0 $X=62830 $Y=318000
X1056 1 2 279 282 280 283 2 275 1 sky130_fd_sc_hd__o22a_4 $T=63020 323680 0 0 $X=62830 $Y=323440
X1057 1 2 290 282 280 288 2 286 1 sky130_fd_sc_hd__o22a_4 $T=72680 323680 0 0 $X=72490 $Y=323440
X1058 1 2 295 282 280 293 2 294 1 sky130_fd_sc_hd__o22a_4 $T=91080 323680 0 0 $X=90890 $Y=323440
X1059 1 2 299 282 280 301 2 292 1 sky130_fd_sc_hd__o22a_4 $T=93840 318240 1 0 $X=93650 $Y=315280
X1060 1 2 304 93 92 302 2 303 1 sky130_fd_sc_hd__o22a_4 $T=115000 318240 1 0 $X=114810 $Y=315280
X1061 1 2 307 93 92 306 2 308 1 sky130_fd_sc_hd__o22a_4 $T=120980 318240 0 0 $X=120790 $Y=318000
X1062 1 2 108 93 109 92 2 312 1 sky130_fd_sc_hd__o22a_4 $T=132940 312800 0 0 $X=132750 $Y=312560
X1063 1 2 115 111 112 117 2 103 1 sky130_fd_sc_hd__o22a_4 $T=139840 312800 1 0 $X=139650 $Y=309840
X1064 1 2 317 111 112 318 2 316 1 sky130_fd_sc_hd__o22a_4 $T=139840 329120 1 0 $X=139650 $Y=326160
X1065 1 2 324 111 112 321 2 319 1 sky130_fd_sc_hd__o22a_4 $T=149960 329120 1 0 $X=149770 $Y=326160
X1066 1 2 325 111 112 323 2 326 1 sky130_fd_sc_hd__o22a_4 $T=156860 318240 0 0 $X=156670 $Y=318000
X1067 1 2 332 111 112 333 2 328 1 sky130_fd_sc_hd__o22a_4 $T=165600 329120 1 0 $X=165410 $Y=326160
X1068 1 2 335 132 131 337 2 336 1 sky130_fd_sc_hd__o22a_4 $T=175260 318240 0 0 $X=175070 $Y=318000
X1069 1 2 340 132 131 343 2 339 1 sky130_fd_sc_hd__o22a_4 $T=185380 318240 0 0 $X=185190 $Y=318000
X1070 1 2 142 150 151 149 2 346 1 sky130_fd_sc_hd__o22a_4 $T=201940 312800 1 0 $X=201750 $Y=309840
X1071 1 2 351 157 159 355 2 354 1 sky130_fd_sc_hd__o22a_4 $T=218500 318240 1 0 $X=218310 $Y=315280
X1072 1 2 357 157 159 356 2 352 1 sky130_fd_sc_hd__o22a_4 $T=222180 329120 1 0 $X=221990 $Y=326160
X1073 1 2 168 157 159 359 2 169 1 sky130_fd_sc_hd__o22a_4 $T=231380 318240 1 0 $X=231190 $Y=315280
X1074 1 2 358 157 159 361 2 362 1 sky130_fd_sc_hd__o22a_4 $T=231380 323680 0 0 $X=231190 $Y=323440
X1075 1 2 370 178 180 369 2 371 1 sky130_fd_sc_hd__o22a_4 $T=253460 318240 1 0 $X=253270 $Y=315280
X1076 1 2 366 178 180 367 2 373 1 sky130_fd_sc_hd__o22a_4 $T=255300 323680 1 0 $X=255110 $Y=320720
X1077 1 2 376 178 180 374 2 375 1 sky130_fd_sc_hd__o22a_4 $T=259440 318240 0 0 $X=259250 $Y=318000
X1078 1 2 213 212 217 208 2 384 1 sky130_fd_sc_hd__o22a_4 $T=303140 312800 1 0 $X=302950 $Y=309840
X1079 1 2 85 2 282 1 sky130_fd_sc_hd__buf_1 $T=105340 312800 1 0 $X=105150 $Y=309840
X1080 1 2 90 2 280 1 sky130_fd_sc_hd__buf_1 $T=109940 312800 1 0 $X=109750 $Y=309840
X1081 1 2 130 2 131 1 sky130_fd_sc_hd__buf_1 $T=175720 312800 1 0 $X=175530 $Y=309840
X1082 1 2 160 2 145 1 sky130_fd_sc_hd__buf_1 $T=219880 312800 1 0 $X=219690 $Y=309840
X1083 1 2 160 2 176 1 sky130_fd_sc_hd__buf_1 $T=273700 312800 1 0 $X=273510 $Y=309840
X1084 1 2 160 2 199 1 sky130_fd_sc_hd__buf_1 $T=284740 312800 1 0 $X=284550 $Y=309840
X1085 1 2 56 279 58 2 283 1 sky130_fd_sc_hd__o21a_4 $T=62100 323680 1 0 $X=61910 $Y=320720
X1086 1 2 57 278 58 2 284 1 sky130_fd_sc_hd__o21a_4 $T=62560 318240 1 0 $X=62370 $Y=315280
X1087 1 2 68 290 58 2 288 1 sky130_fd_sc_hd__o21a_4 $T=77280 323680 1 0 $X=77090 $Y=320720
X1088 1 2 75 295 58 2 293 1 sky130_fd_sc_hd__o21a_4 $T=92920 323680 1 0 $X=92730 $Y=320720
X1089 1 2 89 299 82 2 301 1 sky130_fd_sc_hd__o21a_4 $T=105340 318240 1 0 $X=105150 $Y=315280
X1090 1 2 96 304 82 2 302 1 sky130_fd_sc_hd__o21a_4 $T=119140 312800 0 0 $X=118950 $Y=312560
X1091 1 2 101 307 82 2 306 1 sky130_fd_sc_hd__o21a_4 $T=122360 323680 1 0 $X=122170 $Y=320720
X1092 1 2 56 317 118 2 318 1 sky130_fd_sc_hd__o21a_4 $T=147200 323680 0 0 $X=147010 $Y=323440
X1093 1 2 57 115 118 2 117 1 sky130_fd_sc_hd__o21a_4 $T=149960 312800 1 0 $X=149770 $Y=309840
X1094 1 2 75 324 118 2 321 1 sky130_fd_sc_hd__o21a_4 $T=155480 323680 0 0 $X=155290 $Y=323440
X1095 1 2 68 325 118 2 323 1 sky130_fd_sc_hd__o21a_4 $T=156860 312800 0 0 $X=156670 $Y=312560
X1096 1 2 89 332 129 2 333 1 sky130_fd_sc_hd__o21a_4 $T=173880 323680 1 0 $X=173690 $Y=320720
X1097 1 2 101 335 129 2 337 1 sky130_fd_sc_hd__o21a_4 $T=178940 318240 1 0 $X=178750 $Y=315280
X1098 1 2 139 340 129 2 343 1 sky130_fd_sc_hd__o21a_4 $T=189520 318240 1 0 $X=189330 $Y=315280
X1099 1 2 139 142 148 2 149 1 sky130_fd_sc_hd__o21a_4 $T=203320 312800 0 0 $X=203130 $Y=312560
X1100 1 2 68 351 165 2 355 1 sky130_fd_sc_hd__o21a_4 $T=220800 312800 0 0 $X=220610 $Y=312560
X1101 1 2 57 357 165 2 356 1 sky130_fd_sc_hd__o21a_4 $T=220800 323680 1 0 $X=220610 $Y=320720
X1102 1 2 56 358 165 2 361 1 sky130_fd_sc_hd__o21a_4 $T=230000 323680 1 0 $X=229810 $Y=320720
X1103 1 2 75 168 165 2 359 1 sky130_fd_sc_hd__o21a_4 $T=231840 312800 0 0 $X=231650 $Y=312560
X1104 1 2 175 366 165 2 367 1 sky130_fd_sc_hd__o21a_4 $T=247480 312800 0 0 $X=247290 $Y=312560
X1105 1 2 181 370 183 2 369 1 sky130_fd_sc_hd__o21a_4 $T=253000 312800 1 0 $X=252810 $Y=309840
X1106 1 2 182 376 183 2 374 1 sky130_fd_sc_hd__o21a_4 $T=259440 312800 0 0 $X=259250 $Y=312560
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 4 ICV_7 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3
** N=3 EP=3 IP=9 FDC=3
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 3 sky130_fd_sc_hd__diode_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_24 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249
** N=544 EP=249 IP=6021 FDC=8634
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=265145 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=270585 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=276025 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=281465 $D=191
X4 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=286905 $D=191
X5 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=292345 $D=191
X6 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=297785 $D=191
X7 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=303225 $D=191
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 263840 0 0 $X=5330 $Y=263600
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 296480 1 0 $X=18210 $Y=293520
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 296480 1 0 $X=25570 $Y=293520
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=34040 296480 0 0 $X=33850 $Y=296240
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=46460 280160 1 0 $X=46270 $Y=277200
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=53360 285600 1 0 $X=53170 $Y=282640
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=62100 285600 0 0 $X=61910 $Y=285360
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=68540 280160 1 0 $X=68350 $Y=277200
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=91540 269280 1 0 $X=91350 $Y=266320
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=104420 307360 1 0 $X=104230 $Y=304400
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=132480 296480 1 0 $X=132290 $Y=293520
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 301920 0 0 $X=144250 $Y=301680
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 307360 0 0 $X=144250 $Y=307120
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 280160 1 0 $X=160350 $Y=277200
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=172500 280160 0 0 $X=172310 $Y=279920
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 307360 0 0 $X=174150 $Y=307120
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=197800 291040 1 0 $X=197610 $Y=288080
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=216660 285600 1 0 $X=216470 $Y=282640
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220800 307360 0 0 $X=220610 $Y=307120
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=225400 263840 0 0 $X=225210 $Y=263600
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 274720 1 0 $X=242690 $Y=271760
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=276000 263840 0 0 $X=275810 $Y=263600
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=281520 263840 0 0 $X=281330 $Y=263600
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=283820 301920 1 0 $X=283630 $Y=298960
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286580 307360 0 0 $X=286390 $Y=307120
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=291180 291040 1 0 $X=290990 $Y=288080
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 296480 1 0 $X=314450 $Y=293520
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 296480 0 0 $X=314450 $Y=296240
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 285600 0 0 $X=340670 $Y=285360
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=347760 285600 1 0 $X=347570 $Y=282640
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 263840 1 180 $X=348950 $Y=263600
X39 1 2 ICV_1 $T=5520 269280 1 0 $X=5330 $Y=266320
X40 1 2 ICV_1 $T=5520 274720 1 0 $X=5330 $Y=271760
X41 1 2 ICV_1 $T=5520 280160 1 0 $X=5330 $Y=277200
X42 1 2 ICV_1 $T=5520 285600 1 0 $X=5330 $Y=282640
X43 1 2 ICV_1 $T=5520 291040 1 0 $X=5330 $Y=288080
X44 1 2 ICV_1 $T=5520 296480 1 0 $X=5330 $Y=293520
X45 1 2 ICV_1 $T=5520 301920 1 0 $X=5330 $Y=298960
X46 1 2 ICV_1 $T=5520 307360 1 0 $X=5330 $Y=304400
X47 1 2 ICV_1 $T=6900 307360 1 0 $X=6710 $Y=304400
X48 1 2 ICV_1 $T=350520 269280 0 180 $X=348950 $Y=266320
X49 1 2 ICV_1 $T=350520 274720 0 180 $X=348950 $Y=271760
X50 1 2 ICV_1 $T=350520 280160 0 180 $X=348950 $Y=277200
X51 1 2 ICV_1 $T=350520 285600 0 180 $X=348950 $Y=282640
X52 1 2 ICV_1 $T=350520 291040 0 180 $X=348950 $Y=288080
X53 1 2 ICV_1 $T=350520 296480 0 180 $X=348950 $Y=293520
X54 1 2 ICV_1 $T=350520 301920 0 180 $X=348950 $Y=298960
X55 1 2 ICV_1 $T=350520 307360 0 180 $X=348950 $Y=304400
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 280160 1 0 $X=15910 $Y=277200
X167 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=18400 280160 0 0 $X=18210 $Y=279920
X168 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=27140 263840 0 0 $X=26950 $Y=263600
X169 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 291040 0 0 $X=29710 $Y=290800
X170 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=33120 285600 1 0 $X=32930 $Y=282640
X171 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39100 301920 1 0 $X=38910 $Y=298960
X172 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=41400 291040 1 0 $X=41210 $Y=288080
X173 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=42780 280160 1 0 $X=42590 $Y=277200
X174 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 285600 1 0 $X=43970 $Y=282640
X175 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=45080 274720 0 0 $X=44890 $Y=274480
X176 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=51060 274720 0 0 $X=50870 $Y=274480
X177 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=65780 301920 0 0 $X=65590 $Y=301680
X178 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=70840 291040 0 0 $X=70650 $Y=290800
X179 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 291040 1 0 $X=72030 $Y=288080
X180 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 296480 1 0 $X=72030 $Y=293520
X181 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=75440 280160 0 0 $X=75250 $Y=279920
X182 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=75900 301920 0 0 $X=75710 $Y=301680
X183 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 285600 1 0 $X=76170 $Y=282640
X184 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=77740 307360 0 0 $X=77550 $Y=307120
X185 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=81420 274720 1 0 $X=81230 $Y=271760
X186 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=85560 307360 0 0 $X=85370 $Y=307120
X187 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=87860 269280 1 0 $X=87670 $Y=266320
X188 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=88780 291040 1 0 $X=88590 $Y=288080
X189 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=95680 269280 0 0 $X=95490 $Y=269040
X190 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=95680 280160 0 0 $X=95490 $Y=279920
X191 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=95680 291040 0 0 $X=95490 $Y=290800
X192 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=97060 269280 1 0 $X=96870 $Y=266320
X193 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=97980 291040 1 0 $X=97790 $Y=288080
X194 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=98440 274720 0 0 $X=98250 $Y=274480
X195 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 296480 1 0 $X=100090 $Y=293520
X196 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 307360 1 0 $X=100090 $Y=304400
X197 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 296480 1 0 $X=104230 $Y=293520
X198 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=116380 280160 1 0 $X=116190 $Y=277200
X199 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=116840 274720 1 0 $X=116650 $Y=271760
X200 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=117760 301920 1 0 $X=117570 $Y=298960
X201 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=120980 285600 1 0 $X=120790 $Y=282640
X202 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126960 285600 1 0 $X=126770 $Y=282640
X203 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126960 301920 1 0 $X=126770 $Y=298960
X204 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=135700 269280 0 0 $X=135510 $Y=269040
X205 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=140300 274720 0 0 $X=140110 $Y=274480
X206 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=140760 280160 0 0 $X=140570 $Y=279920
X207 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=140760 301920 0 0 $X=140570 $Y=301680
X208 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142140 296480 0 0 $X=141950 $Y=296240
X209 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=147200 301920 1 0 $X=147010 $Y=298960
X210 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=149960 274720 1 0 $X=149770 $Y=271760
X211 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 269280 1 0 $X=156210 $Y=266320
X212 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=157320 301920 0 0 $X=157130 $Y=301680
X213 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=160540 296480 1 0 $X=160350 $Y=293520
X214 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=164220 301920 0 0 $X=164030 $Y=301680
X215 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 274720 1 0 $X=165410 $Y=271760
X216 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=168820 280160 0 0 $X=168630 $Y=279920
X217 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 263840 0 0 $X=174150 $Y=263600
X218 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178020 285600 1 0 $X=177830 $Y=282640
X219 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=179400 280160 1 0 $X=179210 $Y=277200
X220 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184000 285600 1 0 $X=183810 $Y=282640
X221 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 296480 1 0 $X=184270 $Y=293520
X222 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=185840 296480 0 0 $X=185650 $Y=296240
X223 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 280160 1 0 $X=188410 $Y=277200
X224 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=193660 285600 0 0 $X=193470 $Y=285360
X225 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194120 291040 1 0 $X=193930 $Y=288080
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194580 269280 1 0 $X=194390 $Y=266320
X227 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=200100 301920 1 0 $X=199910 $Y=298960
X228 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211600 280160 1 0 $X=211410 $Y=277200
X229 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 280160 1 0 $X=216470 $Y=277200
X230 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=219420 301920 1 0 $X=219230 $Y=298960
X231 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=219420 307360 1 0 $X=219230 $Y=304400
X232 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=222180 274720 1 0 $X=221990 $Y=271760
X233 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=222180 285600 1 0 $X=221990 $Y=282640
X234 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=225860 301920 1 0 $X=225670 $Y=298960
X235 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 307360 0 0 $X=226130 $Y=307120
X236 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=229540 307360 1 0 $X=229350 $Y=304400
X237 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 280160 0 0 $X=230270 $Y=279920
X238 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 301920 0 0 $X=230270 $Y=301680
X239 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=235520 307360 1 0 $X=235330 $Y=304400
X240 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239200 274720 1 0 $X=239010 $Y=271760
X241 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239660 269280 1 0 $X=239470 $Y=266320
X242 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240120 296480 1 0 $X=239930 $Y=293520
X243 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240120 301920 1 0 $X=239930 $Y=298960
X244 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 307360 1 0 $X=240390 $Y=304400
X245 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=247020 280160 0 0 $X=246830 $Y=279920
X246 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249780 280160 1 0 $X=249590 $Y=277200
X247 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=250240 274720 1 0 $X=250050 $Y=271760
X248 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=253460 263840 0 0 $X=253270 $Y=263600
X249 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254380 280160 0 0 $X=254190 $Y=279920
X250 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=255760 285600 1 0 $X=255570 $Y=282640
X251 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=256220 291040 1 0 $X=256030 $Y=288080
X252 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=264500 291040 0 0 $X=264310 $Y=290800
X253 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267720 296480 1 0 $X=267530 $Y=293520
X254 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 274720 1 0 $X=268450 $Y=271760
X255 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=275080 285600 1 0 $X=274890 $Y=282640
X256 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278300 296480 1 0 $X=278110 $Y=293520
X257 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278760 274720 0 0 $X=278570 $Y=274480
X258 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=279220 269280 1 0 $X=279030 $Y=266320
X259 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=279680 280160 0 0 $X=279490 $Y=279920
X260 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286580 280160 0 0 $X=286390 $Y=279920
X261 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=293480 280160 0 0 $X=293290 $Y=279920
X262 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=294400 301920 1 0 $X=294210 $Y=298960
X263 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=297160 296480 0 0 $X=296970 $Y=296240
X264 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 291040 1 0 $X=300650 $Y=288080
X265 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 280160 0 0 $X=310310 $Y=279920
X266 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310960 291040 1 0 $X=310770 $Y=288080
X267 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 291040 0 0 $X=314450 $Y=290800
X268 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=320160 274720 0 0 $X=319970 $Y=274480
X269 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=323840 274720 1 0 $X=323650 $Y=271760
X270 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=323840 280160 1 0 $X=323650 $Y=277200
X271 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 285600 1 0 $X=328710 $Y=282640
X272 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 291040 1 0 $X=328710 $Y=288080
X273 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 296480 1 0 $X=328710 $Y=293520
X274 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=330740 263840 0 0 $X=330550 $Y=263600
X275 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344080 285600 1 0 $X=343890 $Y=282640
X276 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 269280 1 0 $X=345270 $Y=266320
X277 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 274720 1 0 $X=345270 $Y=271760
X278 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=56120 296480 1 0 $X=55930 $Y=293520
X279 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=60260 285600 1 0 $X=60070 $Y=282640
X280 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=66700 291040 1 0 $X=66510 $Y=288080
X281 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=69920 280160 0 0 $X=69730 $Y=279920
X282 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=70380 301920 1 0 $X=70190 $Y=298960
X283 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=72220 307360 0 0 $X=72030 $Y=307120
X284 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82340 263840 0 0 $X=82150 $Y=263600
X285 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=94760 307360 1 0 $X=94570 $Y=304400
X286 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=114080 307360 1 0 $X=113890 $Y=304400
X287 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=115460 285600 1 0 $X=115270 $Y=282640
X288 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=117760 296480 1 0 $X=117570 $Y=293520
X289 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 280160 1 0 $X=125390 $Y=277200
X290 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=126960 301920 0 0 $X=126770 $Y=301680
X291 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=137540 280160 1 0 $X=137350 $Y=277200
X292 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=141680 301920 1 0 $X=141490 $Y=298960
X293 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=144440 274720 1 0 $X=144250 $Y=271760
X294 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=150880 269280 1 0 $X=150690 $Y=266320
X295 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=151340 263840 0 0 $X=151150 $Y=263600
X296 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=152720 285600 1 0 $X=152530 $Y=282640
X297 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=152720 301920 1 0 $X=152530 $Y=298960
X298 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=153180 296480 1 0 $X=152990 $Y=293520
X299 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=154100 280160 0 0 $X=153910 $Y=279920
X300 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=167900 263840 0 0 $X=167710 $Y=263600
X301 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=180780 291040 1 0 $X=180590 $Y=288080
X302 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=191360 307360 0 0 $X=191170 $Y=307120
X303 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=193660 285600 1 0 $X=193470 $Y=282640
X304 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195500 280160 0 0 $X=195310 $Y=279920
X305 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195960 307360 1 0 $X=195770 $Y=304400
X306 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=207920 301920 1 0 $X=207730 $Y=298960
X307 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210680 274720 1 0 $X=210490 $Y=271760
X308 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210680 307360 1 0 $X=210490 $Y=304400
X309 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=218500 274720 0 0 $X=218310 $Y=274480
X310 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235520 285600 0 0 $X=235330 $Y=285360
X311 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=247940 269280 0 0 $X=247750 $Y=269040
X312 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=247940 296480 0 0 $X=247750 $Y=296240
X313 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=252540 291040 0 0 $X=252350 $Y=290800
X314 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=264040 291040 1 0 $X=263850 $Y=288080
X315 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=265880 285600 1 0 $X=265690 $Y=282640
X316 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=265880 301920 1 0 $X=265690 $Y=298960
X317 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=266340 280160 1 0 $X=266150 $Y=277200
X318 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293940 291040 1 0 $X=293750 $Y=288080
X319 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=320160 285600 1 0 $X=319970 $Y=282640
X320 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=321080 291040 1 0 $X=320890 $Y=288080
X321 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322920 296480 1 0 $X=322730 $Y=293520
X322 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=325220 291040 0 0 $X=325030 $Y=290800
X323 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=327980 269280 0 0 $X=327790 $Y=269040
X324 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=327980 280160 0 0 $X=327790 $Y=279920
X325 1 2 ICV_2 $T=19780 296480 1 0 $X=19590 $Y=293520
X326 1 2 ICV_2 $T=61640 280160 0 0 $X=61450 $Y=279920
X327 1 2 ICV_2 $T=61640 291040 0 0 $X=61450 $Y=290800
X328 1 2 ICV_2 $T=89700 269280 0 0 $X=89510 $Y=269040
X329 1 2 ICV_2 $T=89700 280160 0 0 $X=89510 $Y=279920
X330 1 2 ICV_2 $T=89700 291040 0 0 $X=89510 $Y=290800
X331 1 2 ICV_2 $T=145820 269280 0 0 $X=145630 $Y=269040
X332 1 2 ICV_2 $T=160080 269280 1 0 $X=159890 $Y=266320
X333 1 2 ICV_2 $T=160080 291040 1 0 $X=159890 $Y=288080
X334 1 2 ICV_2 $T=160080 301920 1 0 $X=159890 $Y=298960
X335 1 2 ICV_2 $T=188140 291040 1 0 $X=187950 $Y=288080
X336 1 2 ICV_2 $T=216200 274720 1 0 $X=216010 $Y=271760
X337 1 2 ICV_2 $T=244260 269280 1 0 $X=244070 $Y=266320
X338 1 2 ICV_2 $T=244260 274720 1 0 $X=244070 $Y=271760
X339 1 2 ICV_2 $T=244260 301920 1 0 $X=244070 $Y=298960
X340 1 2 ICV_2 $T=244260 307360 1 0 $X=244070 $Y=304400
X341 1 2 ICV_2 $T=272320 296480 1 0 $X=272130 $Y=293520
X342 1 2 ICV_2 $T=272320 301920 1 0 $X=272130 $Y=298960
X343 1 2 ICV_2 $T=314180 274720 0 0 $X=313990 $Y=274480
X344 1 2 ICV_2 $T=328440 269280 1 0 $X=328250 $Y=266320
X345 1 2 ICV_2 $T=342240 263840 0 0 $X=342050 $Y=263600
X346 1 2 ICV_2 $T=342240 269280 0 0 $X=342050 $Y=269040
X347 1 2 ICV_2 $T=342240 274720 0 0 $X=342050 $Y=274480
X348 1 2 ICV_2 $T=342240 280160 0 0 $X=342050 $Y=279920
X349 1 2 ICV_2 $T=342240 285600 0 0 $X=342050 $Y=285360
X350 1 2 ICV_2 $T=342240 291040 0 0 $X=342050 $Y=290800
X351 1 2 ICV_2 $T=342240 296480 0 0 $X=342050 $Y=296240
X352 1 2 ICV_2 $T=342240 307360 0 0 $X=342050 $Y=307120
X353 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=10580 269280 1 0 $X=10390 $Y=266320
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 274720 1 0 $X=17750 $Y=271760
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 285600 1 0 $X=17750 $Y=282640
X356 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 301920 1 0 $X=17750 $Y=298960
X357 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 269280 0 0 $X=18210 $Y=269040
X358 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 274720 0 0 $X=18210 $Y=274480
X359 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31280 285600 0 0 $X=31090 $Y=285360
X360 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31280 301920 0 0 $X=31090 $Y=301680
X361 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 280160 1 0 $X=31550 $Y=277200
X362 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=37260 274720 1 0 $X=37070 $Y=271760
X363 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=37260 307360 1 0 $X=37070 $Y=304400
X364 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=38180 269280 1 0 $X=37990 $Y=266320
X365 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=45540 263840 0 0 $X=45350 $Y=263600
X366 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 296480 1 0 $X=45810 $Y=293520
X367 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=55660 269280 0 0 $X=55470 $Y=269040
X368 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=57500 301920 0 0 $X=57310 $Y=301680
X369 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59340 263840 0 0 $X=59150 $Y=263600
X370 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=61640 296480 1 0 $X=61450 $Y=293520
X371 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=63020 291040 1 0 $X=62830 $Y=288080
X372 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69920 269280 1 0 $X=69730 $Y=266320
X373 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=72220 263840 0 0 $X=72030 $Y=263600
X374 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87860 263840 0 0 $X=87670 $Y=263600
X375 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=97980 307360 0 0 $X=97790 $Y=307120
X376 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 280160 1 0 $X=101930 $Y=277200
X377 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104880 285600 0 0 $X=104690 $Y=285360
X378 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=106720 301920 1 0 $X=106530 $Y=298960
X379 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=108100 280160 0 0 $X=107910 $Y=279920
X380 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=112700 263840 0 0 $X=112510 $Y=263600
X381 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 274720 0 0 $X=115730 $Y=274480
X382 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=132480 291040 1 0 $X=132290 $Y=288080
X383 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=132480 301920 0 0 $X=132290 $Y=301680
X384 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=135700 307360 0 0 $X=135510 $Y=307120
X385 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=150880 307360 0 0 $X=150690 $Y=307120
X386 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=156860 263840 0 0 $X=156670 $Y=263600
X387 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 285600 1 0 $X=158050 $Y=282640
X388 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 301920 1 0 $X=158050 $Y=298960
X389 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 307360 1 0 $X=158050 $Y=304400
X390 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=166060 291040 1 0 $X=165870 $Y=288080
X391 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 307360 1 0 $X=171850 $Y=304400
X392 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=184460 269280 0 0 $X=184270 $Y=269040
X393 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 291040 1 0 $X=186110 $Y=288080
X394 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186760 280160 0 0 $X=186570 $Y=279920
X395 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=197800 296480 0 0 $X=197610 $Y=296240
X396 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=211600 291040 0 0 $X=211410 $Y=290800
X397 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=213440 280160 0 0 $X=213250 $Y=279920
X398 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=218960 269280 1 0 $X=218770 $Y=266320
X399 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=224020 291040 0 0 $X=223830 $Y=290800
X400 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=227700 301920 0 0 $X=227510 $Y=301680
X401 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230460 296480 0 0 $X=230270 $Y=296240
X402 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=234600 280160 1 0 $X=234410 $Y=277200
X403 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=241960 285600 1 0 $X=241770 $Y=282640
X404 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244260 291040 0 0 $X=244070 $Y=290800
X405 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=252540 285600 0 0 $X=252350 $Y=285360
X406 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258060 301920 1 0 $X=257870 $Y=298960
X407 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=264960 269280 1 0 $X=264770 $Y=266320
X408 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=270020 269280 1 0 $X=269830 $Y=266320
X409 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284280 291040 1 0 $X=284090 $Y=288080
X410 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=285660 280160 1 0 $X=285470 $Y=277200
X411 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=287500 274720 1 0 $X=287310 $Y=271760
X412 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=289340 269280 1 0 $X=289150 $Y=266320
X413 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=289340 307360 1 0 $X=289150 $Y=304400
X414 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=296240 280160 1 0 $X=296050 $Y=277200
X415 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 285600 1 0 $X=298350 $Y=282640
X416 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=303600 285600 0 0 $X=303410 $Y=285360
X417 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=304520 280160 1 0 $X=304330 $Y=277200
X418 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=310040 269280 0 0 $X=309850 $Y=269040
X419 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=314640 269280 0 0 $X=314450 $Y=269040
X420 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 269280 1 0 $X=325950 $Y=266320
X421 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 291040 1 0 $X=326410 $Y=288080
X422 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 301920 1 0 $X=326410 $Y=298960
X423 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 307360 1 0 $X=328710 $Y=304400
X424 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=330740 291040 0 0 $X=330550 $Y=290800
X425 1 3 sky130_fd_sc_hd__diode_2 $T=7820 285600 0 0 $X=7630 $Y=285360
X426 1 3 sky130_fd_sc_hd__diode_2 $T=11040 263840 0 0 $X=10850 $Y=263600
X427 1 5 sky130_fd_sc_hd__diode_2 $T=36340 291040 0 0 $X=36150 $Y=290800
X428 1 32 sky130_fd_sc_hd__diode_2 $T=37260 269280 0 0 $X=37070 $Y=269040
X429 1 330 sky130_fd_sc_hd__diode_2 $T=46460 285600 0 0 $X=46270 $Y=285360
X430 1 40 sky130_fd_sc_hd__diode_2 $T=48300 269280 0 0 $X=48110 $Y=269040
X431 1 336 sky130_fd_sc_hd__diode_2 $T=50600 280160 1 0 $X=50410 $Y=277200
X432 1 336 sky130_fd_sc_hd__diode_2 $T=56580 274720 1 0 $X=56390 $Y=271760
X433 1 34 sky130_fd_sc_hd__diode_2 $T=56580 307360 1 0 $X=56390 $Y=304400
X434 1 50 sky130_fd_sc_hd__diode_2 $T=57960 280160 0 0 $X=57770 $Y=279920
X435 1 5 sky130_fd_sc_hd__diode_2 $T=63940 296480 1 0 $X=63750 $Y=293520
X436 1 319 sky130_fd_sc_hd__diode_2 $T=69920 301920 0 0 $X=69730 $Y=301680
X437 1 63 sky130_fd_sc_hd__diode_2 $T=70380 269280 0 0 $X=70190 $Y=269040
X438 1 336 sky130_fd_sc_hd__diode_2 $T=72220 280160 1 0 $X=72030 $Y=277200
X439 1 351 sky130_fd_sc_hd__diode_2 $T=75440 291040 0 0 $X=75250 $Y=290800
X440 1 360 sky130_fd_sc_hd__diode_2 $T=78660 301920 1 0 $X=78470 $Y=298960
X441 1 42 sky130_fd_sc_hd__diode_2 $T=81880 269280 0 0 $X=81690 $Y=269040
X442 1 357 sky130_fd_sc_hd__diode_2 $T=86020 291040 0 0 $X=85830 $Y=290800
X443 1 5 sky130_fd_sc_hd__diode_2 $T=99820 291040 0 0 $X=99630 $Y=290800
X444 1 76 sky130_fd_sc_hd__diode_2 $T=101660 285600 0 0 $X=101470 $Y=285360
X445 1 74 sky130_fd_sc_hd__diode_2 $T=102580 301920 0 0 $X=102390 $Y=301680
X446 1 78 sky130_fd_sc_hd__diode_2 $T=103960 307360 0 0 $X=103770 $Y=307120
X447 1 377 sky130_fd_sc_hd__diode_2 $T=104420 269280 0 0 $X=104230 $Y=269040
X448 1 382 sky130_fd_sc_hd__diode_2 $T=123740 274720 0 0 $X=123550 $Y=274480
X449 1 5 sky130_fd_sc_hd__diode_2 $T=124200 285600 0 0 $X=124010 $Y=285360
X450 1 384 sky130_fd_sc_hd__diode_2 $T=124660 263840 0 0 $X=124470 $Y=263600
X451 1 5 sky130_fd_sc_hd__diode_2 $T=124660 291040 0 0 $X=124470 $Y=290800
X452 1 5 sky130_fd_sc_hd__diode_2 $T=127880 274720 0 0 $X=127690 $Y=274480
X453 1 359 sky130_fd_sc_hd__diode_2 $T=141680 291040 0 0 $X=141490 $Y=290800
X454 1 5 sky130_fd_sc_hd__diode_2 $T=151800 274720 0 0 $X=151610 $Y=274480
X455 1 114 sky130_fd_sc_hd__diode_2 $T=153640 291040 0 0 $X=153450 $Y=290800
X456 1 115 sky130_fd_sc_hd__diode_2 $T=160540 307360 0 0 $X=160350 $Y=307120
X457 1 405 sky130_fd_sc_hd__diode_2 $T=164220 269280 0 0 $X=164030 $Y=269040
X458 1 125 sky130_fd_sc_hd__diode_2 $T=164220 307360 0 0 $X=164030 $Y=307120
X459 1 123 sky130_fd_sc_hd__diode_2 $T=166060 269280 1 0 $X=165870 $Y=266320
X460 1 120 sky130_fd_sc_hd__diode_2 $T=177560 285600 0 0 $X=177370 $Y=285360
X461 1 5 sky130_fd_sc_hd__diode_2 $T=181240 285600 0 0 $X=181050 $Y=285360
X462 1 415 sky130_fd_sc_hd__diode_2 $T=182160 301920 1 0 $X=181970 $Y=298960
X463 1 139 sky130_fd_sc_hd__diode_2 $T=186760 269280 0 0 $X=186570 $Y=269040
X464 1 80 sky130_fd_sc_hd__diode_2 $T=187680 301920 0 0 $X=187490 $Y=301680
X465 1 423 sky130_fd_sc_hd__diode_2 $T=196880 274720 1 0 $X=196690 $Y=271760
X466 1 145 sky130_fd_sc_hd__diode_2 $T=199180 285600 1 0 $X=198990 $Y=282640
X467 1 425 sky130_fd_sc_hd__diode_2 $T=200560 296480 1 0 $X=200370 $Y=293520
X468 1 80 sky130_fd_sc_hd__diode_2 $T=203320 291040 0 0 $X=203130 $Y=290800
X469 1 150 sky130_fd_sc_hd__diode_2 $T=205160 274720 1 0 $X=204970 $Y=271760
X470 1 152 sky130_fd_sc_hd__diode_2 $T=219420 280160 0 0 $X=219230 $Y=279920
X471 1 444 sky130_fd_sc_hd__diode_2 $T=226320 291040 0 0 $X=226130 $Y=290800
X472 1 5 sky130_fd_sc_hd__diode_2 $T=234600 280160 0 0 $X=234410 $Y=279920
X473 1 5 sky130_fd_sc_hd__diode_2 $T=236900 263840 0 0 $X=236710 $Y=263600
X474 1 124 sky130_fd_sc_hd__diode_2 $T=238280 291040 0 0 $X=238090 $Y=290800
X475 1 172 sky130_fd_sc_hd__diode_2 $T=248400 307360 0 0 $X=248210 $Y=307120
X476 1 464 sky130_fd_sc_hd__diode_2 $T=262200 263840 0 0 $X=262010 $Y=263600
X477 1 181 sky130_fd_sc_hd__diode_2 $T=265880 301920 0 0 $X=265690 $Y=301680
X478 1 130 sky130_fd_sc_hd__diode_2 $T=266340 263840 0 0 $X=266150 $Y=263600
X479 1 192 sky130_fd_sc_hd__diode_2 $T=272780 274720 0 0 $X=272590 $Y=274480
X480 1 469 sky130_fd_sc_hd__diode_2 $T=273700 274720 1 0 $X=273510 $Y=271760
X481 1 474 sky130_fd_sc_hd__diode_2 $T=281060 307360 1 0 $X=280870 $Y=304400
X482 1 160 sky130_fd_sc_hd__diode_2 $T=287500 296480 0 0 $X=287310 $Y=296240
X483 1 479 sky130_fd_sc_hd__diode_2 $T=287960 280160 1 0 $X=287770 $Y=277200
X484 1 144 sky130_fd_sc_hd__diode_2 $T=288880 274720 0 0 $X=288690 $Y=274480
X485 1 200 sky130_fd_sc_hd__diode_2 $T=293940 285600 0 0 $X=293750 $Y=285360
X486 1 426 sky130_fd_sc_hd__diode_2 $T=298080 285600 0 0 $X=297890 $Y=285360
X487 1 216 sky130_fd_sc_hd__diode_2 $T=300840 301920 0 0 $X=300650 $Y=301680
X488 1 209 sky130_fd_sc_hd__diode_2 $T=304520 296480 0 0 $X=304330 $Y=296240
X489 1 485 sky130_fd_sc_hd__diode_2 $T=308200 301920 1 0 $X=308010 $Y=298960
X490 1 5 sky130_fd_sc_hd__diode_2 $T=331200 307360 1 0 $X=331010 $Y=304400
X491 1 237 sky130_fd_sc_hd__diode_2 $T=338560 263840 0 0 $X=338370 $Y=263600
X492 1 238 sky130_fd_sc_hd__diode_2 $T=338560 269280 0 0 $X=338370 $Y=269040
X493 1 2 4 ICV_4 $T=7820 263840 0 0 $X=7630 $Y=263600
X494 1 2 326 ICV_4 $T=37260 285600 1 0 $X=37070 $Y=282640
X495 1 2 41 ICV_4 $T=49220 301920 1 0 $X=49030 $Y=298960
X496 1 2 47 ICV_4 $T=52900 269280 1 0 $X=52710 $Y=266320
X497 1 2 48 ICV_4 $T=58880 291040 0 0 $X=58690 $Y=290800
X498 1 2 347 ICV_4 $T=60720 301920 1 0 $X=60530 $Y=298960
X499 1 2 354 ICV_4 $T=74980 274720 0 0 $X=74790 $Y=274480
X500 1 2 64 ICV_4 $T=78660 269280 0 0 $X=78470 $Y=269040
X501 1 2 64 ICV_4 $T=91080 274720 0 0 $X=90890 $Y=274480
X502 1 2 82 ICV_4 $T=105800 307360 1 0 $X=105610 $Y=304400
X503 1 2 84 ICV_4 $T=106720 280160 1 0 $X=106530 $Y=277200
X504 1 2 55 ICV_4 $T=108560 269280 0 0 $X=108370 $Y=269040
X505 1 2 379 ICV_4 $T=108560 301920 1 0 $X=108370 $Y=298960
X506 1 2 382 ICV_4 $T=112700 274720 1 0 $X=112510 $Y=271760
X507 1 2 317 ICV_4 $T=113160 291040 0 0 $X=112970 $Y=290800
X508 1 2 381 ICV_4 $T=113160 296480 1 0 $X=112970 $Y=293520
X509 1 2 377 ICV_4 $T=114540 263840 0 0 $X=114350 $Y=263600
X510 1 2 76 ICV_4 $T=121440 291040 0 0 $X=121250 $Y=290800
X511 1 2 381 ICV_4 $T=125120 296480 0 0 $X=124930 $Y=296240
X512 1 2 393 ICV_4 $T=133400 301920 1 0 $X=133210 $Y=298960
X513 1 2 390 ICV_4 $T=138920 296480 1 0 $X=138730 $Y=293520
X514 1 2 394 ICV_4 $T=147200 285600 0 0 $X=147010 $Y=285360
X515 1 2 396 ICV_4 $T=149040 296480 1 0 $X=148850 $Y=293520
X516 1 2 114 ICV_4 $T=155480 307360 0 0 $X=155290 $Y=307120
X517 1 2 399 ICV_4 $T=157780 291040 0 0 $X=157590 $Y=290800
X518 1 2 406 ICV_4 $T=171120 269280 0 0 $X=170930 $Y=269040
X519 1 2 114 ICV_4 $T=171120 274720 0 0 $X=170930 $Y=274480
X520 1 2 399 ICV_4 $T=171120 301920 0 0 $X=170930 $Y=301680
X521 1 2 410 ICV_4 $T=176640 296480 1 0 $X=176450 $Y=293520
X522 1 2 127 ICV_4 $T=177560 307360 1 0 $X=177370 $Y=304400
X523 1 2 409 ICV_4 $T=178940 269280 1 0 $X=178750 $Y=266320
X524 1 2 402 ICV_4 $T=183540 274720 1 0 $X=183350 $Y=271760
X525 1 2 121 ICV_4 $T=189520 263840 0 0 $X=189330 $Y=263600
X526 1 2 134 ICV_4 $T=198720 269280 1 0 $X=198530 $Y=266320
X527 1 2 144 ICV_4 $T=198720 269280 0 0 $X=198530 $Y=269040
X528 1 2 5 ICV_4 $T=198720 274720 0 0 $X=198530 $Y=274480
X529 1 2 148 ICV_4 $T=201940 307360 1 0 $X=201750 $Y=304400
X530 1 2 146 ICV_4 $T=209300 296480 0 0 $X=209110 $Y=296240
X531 1 2 158 ICV_4 $T=213440 269280 1 0 $X=213250 $Y=266320
X532 1 2 120 ICV_4 $T=214820 296480 0 0 $X=214630 $Y=296240
X533 1 2 435 ICV_4 $T=217580 296480 0 0 $X=217390 $Y=296240
X534 1 2 438 ICV_4 $T=221260 280160 1 0 $X=221070 $Y=277200
X535 1 2 5 ICV_4 $T=226780 263840 0 0 $X=226590 $Y=263600
X536 1 2 444 ICV_4 $T=234140 301920 0 0 $X=233950 $Y=301680
X537 1 2 453 ICV_4 $T=250240 307360 1 0 $X=250050 $Y=304400
X538 1 2 459 ICV_4 $T=255300 274720 0 0 $X=255110 $Y=274480
X539 1 2 58 ICV_4 $T=255300 307360 0 0 $X=255110 $Y=307120
X540 1 2 185 ICV_4 $T=259440 263840 0 0 $X=259250 $Y=263600
X541 1 2 46 ICV_4 $T=260360 296480 1 0 $X=260170 $Y=293520
X542 1 2 458 ICV_4 $T=266340 307360 1 0 $X=266150 $Y=304400
X543 1 2 191 ICV_4 $T=269100 307360 1 0 $X=268910 $Y=304400
X544 1 2 445 ICV_4 $T=270020 301920 0 0 $X=269830 $Y=301680
X545 1 2 318 ICV_4 $T=281060 285600 1 0 $X=280870 $Y=282640
X546 1 2 462 ICV_4 $T=282900 263840 0 0 $X=282710 $Y=263600
X547 1 2 159 ICV_4 $T=282900 301920 0 0 $X=282710 $Y=301680
X548 1 2 462 ICV_4 $T=289800 274720 1 0 $X=289610 $Y=271760
X549 1 2 192 ICV_4 $T=293020 307360 0 0 $X=292830 $Y=307120
X550 1 2 192 ICV_4 $T=293940 269280 0 0 $X=293750 $Y=269040
X551 1 2 186 ICV_4 $T=297160 274720 0 0 $X=296970 $Y=274480
X552 1 2 485 ICV_4 $T=301760 269280 1 0 $X=301570 $Y=266320
X553 1 2 489 ICV_4 $T=309120 285600 0 0 $X=308930 $Y=285360
X554 1 2 210 ICV_4 $T=310960 274720 0 0 $X=310770 $Y=274480
X555 1 2 5 ICV_4 $T=311420 263840 0 0 $X=311230 $Y=263600
X556 1 2 225 ICV_4 $T=311420 296480 0 0 $X=311230 $Y=296240
X557 1 2 5 ICV_4 $T=316020 296480 1 0 $X=315830 $Y=293520
X558 1 2 3 ICV_4 $T=332120 274720 1 0 $X=331930 $Y=271760
X559 1 2 5 ICV_4 $T=339480 274720 0 0 $X=339290 $Y=274480
X560 1 2 3 ICV_4 $T=339480 301920 0 0 $X=339290 $Y=301680
X561 1 2 3 ICV_4 $T=339480 307360 0 0 $X=339290 $Y=307120
X562 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 291040 1 0 $X=6710 $Y=288080
X563 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 296480 1 0 $X=6710 $Y=293520
X564 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=18400 301920 0 0 $X=18210 $Y=301680
X565 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30360 274720 0 0 $X=30170 $Y=274480
X566 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30360 307360 0 0 $X=30170 $Y=307120
X567 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30820 269280 0 0 $X=30630 $Y=269040
X568 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=34040 269280 0 0 $X=33850 $Y=269040
X569 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=36340 301920 0 0 $X=36150 $Y=301680
X570 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=41860 301920 0 0 $X=41670 $Y=301680
X571 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=51520 280160 1 0 $X=51330 $Y=277200
X572 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58880 280160 0 0 $X=58690 $Y=279920
X573 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58880 296480 0 0 $X=58690 $Y=296240
X574 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=64860 296480 1 0 $X=64670 $Y=293520
X575 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=65780 285600 1 0 $X=65590 $Y=282640
X576 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 280160 1 0 $X=72950 $Y=277200
X577 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 285600 1 0 $X=72950 $Y=282640
X578 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=86480 280160 0 0 $X=86290 $Y=279920
X579 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=86940 291040 0 0 $X=86750 $Y=290800
X580 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=87400 280160 1 0 $X=87210 $Y=277200
X581 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=87400 307360 1 0 $X=87210 $Y=304400
X582 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101200 274720 1 0 $X=101010 $Y=271760
X583 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101200 301920 1 0 $X=101010 $Y=298960
X584 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=111780 269280 1 0 $X=111590 $Y=266320
X585 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=124660 274720 0 0 $X=124470 $Y=274480
X586 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129260 280160 0 0 $X=129070 $Y=279920
X587 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=161460 307360 0 0 $X=161270 $Y=307120
X588 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=165140 285600 0 0 $X=164950 $Y=285360
X589 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=166980 269280 1 0 $X=166790 $Y=266320
X590 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=173420 285600 1 0 $X=173230 $Y=282640
X591 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=176180 274720 1 0 $X=175990 $Y=271760
X592 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=178480 285600 0 0 $X=178290 $Y=285360
X593 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=183080 301920 1 0 $X=182890 $Y=298960
X594 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=198720 301920 0 0 $X=198530 $Y=301680
X595 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 301920 0 0 $X=202210 $Y=301680
X596 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=206080 274720 1 0 $X=205890 $Y=271760
X597 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=211140 291040 1 0 $X=210950 $Y=288080
X598 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=211600 285600 1 0 $X=211410 $Y=282640
X599 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213440 301920 1 0 $X=213250 $Y=298960
X600 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=223100 296480 1 0 $X=222910 $Y=293520
X601 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 269280 0 0 $X=226590 $Y=269040
X602 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 274720 0 0 $X=226590 $Y=274480
X603 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=227240 291040 0 0 $X=227050 $Y=290800
X604 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=230000 274720 1 0 $X=229810 $Y=271760
X605 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241040 291040 1 0 $X=240850 $Y=288080
X606 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241500 274720 0 0 $X=241310 $Y=274480
X607 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=263120 263840 0 0 $X=262930 $Y=263600
X608 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269560 274720 0 0 $X=269370 $Y=274480
X609 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269560 280160 0 0 $X=269370 $Y=279920
X610 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269560 291040 1 0 $X=269370 $Y=288080
X611 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=277840 307360 1 0 $X=277650 $Y=304400
X612 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=278300 301920 1 0 $X=278110 $Y=298960
X613 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=279680 307360 0 0 $X=279490 $Y=307120
X614 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=281060 280160 1 0 $X=280870 $Y=277200
X615 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=281980 274720 1 0 $X=281790 $Y=271760
X616 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=288420 296480 1 0 $X=288230 $Y=293520
X617 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=293940 307360 1 0 $X=293750 $Y=304400
X618 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=313260 285600 1 0 $X=313070 $Y=282640
X619 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325680 285600 1 0 $X=325490 $Y=282640
X620 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 263840 0 0 $X=339290 $Y=263600
X621 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 269280 0 0 $X=339290 $Y=269040
X622 1 2 322 ICV_6 $T=26220 280160 0 0 $X=26030 $Y=279920
X623 1 2 325 ICV_6 $T=34040 280160 1 0 $X=33850 $Y=277200
X624 1 2 327 ICV_6 $T=38640 296480 1 0 $X=38450 $Y=293520
X625 1 2 328 ICV_6 $T=43240 301920 1 0 $X=43050 $Y=298960
X626 1 2 358 ICV_6 $T=77280 291040 1 0 $X=77090 $Y=288080
X627 1 2 363 ICV_6 $T=96140 285600 0 0 $X=95950 $Y=285360
X628 1 2 370 ICV_6 $T=98440 296480 0 0 $X=98250 $Y=296240
X629 1 2 86 ICV_6 $T=113160 301920 0 0 $X=112970 $Y=301680
X630 1 2 88 ICV_6 $T=113160 307360 0 0 $X=112970 $Y=307120
X631 1 2 92 ICV_6 $T=119140 263840 0 0 $X=118950 $Y=263600
X632 1 2 385 ICV_6 $T=121900 269280 1 0 $X=121710 $Y=266320
X633 1 2 97 ICV_6 $T=126500 269280 1 0 $X=126310 $Y=266320
X634 1 2 95 ICV_6 $T=126960 307360 1 0 $X=126770 $Y=304400
X635 1 2 102 ICV_6 $T=137540 285600 0 0 $X=137350 $Y=285360
X636 1 2 103 ICV_6 $T=140300 269280 0 0 $X=140110 $Y=269040
X637 1 2 397 ICV_6 $T=147200 274720 0 0 $X=147010 $Y=274480
X638 1 2 364 ICV_6 $T=147200 296480 0 0 $X=147010 $Y=296240
X639 1 2 400 ICV_6 $T=153640 274720 1 0 $X=153450 $Y=271760
X640 1 2 407 ICV_6 $T=166980 291040 0 0 $X=166790 $Y=290800
X641 1 2 120 ICV_6 $T=168360 285600 0 0 $X=168170 $Y=285360
X642 1 2 134 ICV_6 $T=178940 274720 1 0 $X=178750 $Y=271760
X643 1 2 418 ICV_6 $T=183540 280160 1 0 $X=183350 $Y=277200
X644 1 2 151 ICV_6 $T=208840 296480 1 0 $X=208650 $Y=293520
X645 1 2 164 ICV_6 $T=221260 269280 1 0 $X=221070 $Y=266320
X646 1 2 151 ICV_6 $T=222180 285600 0 0 $X=221990 $Y=285360
X647 1 2 162 ICV_6 $T=222640 296480 0 0 $X=222450 $Y=296240
X648 1 2 441 ICV_6 $T=231380 263840 0 0 $X=231190 $Y=263600
X649 1 2 173 ICV_6 $T=235520 307360 0 0 $X=235330 $Y=307120
X650 1 2 159 ICV_6 $T=243340 307360 0 0 $X=243150 $Y=307120
X651 1 2 445 ICV_6 $T=272780 280160 0 0 $X=272590 $Y=279920
X652 1 2 468 ICV_6 $T=272780 301920 0 0 $X=272590 $Y=301680
X653 1 2 475 ICV_6 $T=286580 291040 1 0 $X=286390 $Y=288080
X654 1 2 491 ICV_6 $T=308200 274720 1 0 $X=308010 $Y=271760
X655 1 2 472 ICV_6 $T=308200 291040 0 0 $X=308010 $Y=290800
X656 1 2 468 ICV_6 $T=336260 285600 0 0 $X=336070 $Y=285360
X657 1 2 501 ICV_6 $T=336720 291040 0 0 $X=336530 $Y=290800
X658 1 2 446 ICV_6 $T=337180 280160 0 0 $X=336990 $Y=279920
X659 1 2 236 ICV_6 $T=343620 301920 0 0 $X=343430 $Y=301680
X660 1 3 5 ICV_7 $T=7820 269280 1 0 $X=7630 $Y=266320
X661 1 3 5 ICV_7 $T=7820 274720 1 0 $X=7630 $Y=271760
X662 1 5 5 ICV_7 $T=7820 285600 1 0 $X=7630 $Y=282640
X663 1 3 5 ICV_7 $T=7820 301920 1 0 $X=7630 $Y=298960
X664 1 3 5 ICV_7 $T=8280 307360 1 0 $X=8090 $Y=304400
X665 1 3 5 ICV_7 $T=20240 274720 0 0 $X=20050 $Y=274480
X666 1 3 5 ICV_7 $T=20700 269280 0 0 $X=20510 $Y=269040
X667 1 3 5 ICV_7 $T=21160 285600 0 0 $X=20970 $Y=285360
X668 1 3 5 ICV_7 $T=21160 301920 0 0 $X=20970 $Y=301680
X669 1 3 5 ICV_7 $T=22540 280160 0 0 $X=22350 $Y=279920
X670 1 3 5 ICV_7 $T=24380 263840 0 0 $X=24190 $Y=263600
X671 1 5 323 ICV_7 $T=27140 291040 0 0 $X=26950 $Y=290800
X672 1 29 33 ICV_7 $T=34960 307360 0 0 $X=34770 $Y=307120
X673 1 34 330 ICV_7 $T=38640 307360 0 0 $X=38450 $Y=307120
X674 1 29 332 ICV_7 $T=39100 301920 0 0 $X=38910 $Y=301680
X675 1 22 331 ICV_7 $T=42780 285600 0 0 $X=42590 $Y=285360
X676 1 37 338 ICV_7 $T=43240 296480 1 0 $X=43050 $Y=293520
X677 1 335 38 ICV_7 $T=44160 307360 1 0 $X=43970 $Y=304400
X678 1 337 37 ICV_7 $T=44620 301920 0 0 $X=44430 $Y=301680
X679 1 342 42 ICV_7 $T=47840 263840 0 0 $X=47650 $Y=263600
X680 1 330 43 ICV_7 $T=48300 301920 0 0 $X=48110 $Y=301680
X681 1 343 37 ICV_7 $T=50600 285600 1 0 $X=50410 $Y=282640
X682 1 47 343 ICV_7 $T=54740 280160 1 0 $X=54550 $Y=277200
X683 1 5 345 ICV_7 $T=56580 263840 0 0 $X=56390 $Y=263600
X684 1 340 340 ICV_7 $T=57960 269280 0 0 $X=57770 $Y=269040
X685 1 330 37 ICV_7 $T=63020 301920 0 0 $X=62830 $Y=301680
X686 1 56 58 ICV_7 $T=63020 307360 0 0 $X=62830 $Y=307120
X687 1 336 340 ICV_7 $T=65780 274720 1 0 $X=65590 $Y=271760
X688 1 57 55 ICV_7 $T=65780 285600 0 0 $X=65590 $Y=285360
X689 1 49 61 ICV_7 $T=67160 269280 1 0 $X=66970 $Y=266320
X690 1 351 353 ICV_7 $T=68080 291040 0 0 $X=67890 $Y=290800
X691 1 59 61 ICV_7 $T=69460 263840 0 0 $X=69270 $Y=263600
X692 1 350 352 ICV_7 $T=72220 269280 1 0 $X=72030 $Y=266320
X693 1 356 5 ICV_7 $T=74520 263840 0 0 $X=74330 $Y=263600
X694 1 58 364 ICV_7 $T=82340 291040 0 0 $X=82150 $Y=290800
X695 1 359 361 ICV_7 $T=83720 285600 0 0 $X=83530 $Y=285360
X696 1 5 366 ICV_7 $T=86020 269280 0 0 $X=85830 $Y=269040
X697 1 367 5 ICV_7 $T=86020 301920 0 0 $X=85830 $Y=301680
X698 1 371 64 ICV_7 $T=91080 263840 0 0 $X=90890 $Y=263600
X699 1 48 364 ICV_7 $T=92460 285600 0 0 $X=92270 $Y=285360
X700 1 73 75 ICV_7 $T=99820 263840 0 0 $X=99630 $Y=263600
X701 1 373 64 ICV_7 $T=100280 280160 0 0 $X=100090 $Y=279920
X702 1 374 77 ICV_7 $T=100280 307360 0 0 $X=100090 $Y=307120
X703 1 372 80 ICV_7 $T=103040 274720 0 0 $X=102850 $Y=274480
X704 1 377 81 ICV_7 $T=103500 263840 0 0 $X=103310 $Y=263600
X705 1 81 87 ICV_7 $T=109480 301920 0 0 $X=109290 $Y=301680
X706 1 377 75 ICV_7 $T=113160 274720 0 0 $X=112970 $Y=274480
X707 1 57 62 ICV_7 $T=113620 269280 0 0 $X=113430 $Y=269040
X708 1 78 82 ICV_7 $T=113620 296480 0 0 $X=113430 $Y=296240
X709 1 93 84 ICV_7 $T=120060 274720 0 0 $X=119870 $Y=274480
X710 1 80 87 ICV_7 $T=121440 296480 0 0 $X=121250 $Y=296240
X711 1 77 5 ICV_7 $T=121440 307360 0 0 $X=121250 $Y=307120
X712 1 390 359 ICV_7 $T=128340 296480 0 0 $X=128150 $Y=296240
X713 1 95 361 ICV_7 $T=138000 291040 0 0 $X=137810 $Y=290800
X714 1 105 107 ICV_7 $T=138000 307360 0 0 $X=137810 $Y=307120
X715 1 44 106 ICV_7 $T=139380 296480 0 0 $X=139190 $Y=296240
X716 1 108 104 ICV_7 $T=141680 307360 0 0 $X=141490 $Y=307120
X717 1 111 112 ICV_7 $T=148120 301920 0 0 $X=147930 $Y=301680
X718 1 106 50 ICV_7 $T=148120 307360 0 0 $X=147930 $Y=307120
X719 1 121 122 ICV_7 $T=159620 280160 0 0 $X=159430 $Y=279920
X720 1 5 404 ICV_7 $T=161460 301920 0 0 $X=161270 $Y=301680
X721 1 121 5 ICV_7 $T=163300 291040 0 0 $X=163110 $Y=290800
X722 1 406 401 ICV_7 $T=165140 274720 0 0 $X=164950 $Y=274480
X723 1 408 114 ICV_7 $T=166060 301920 1 0 $X=165870 $Y=298960
X724 1 128 115 ICV_7 $T=173880 307360 1 0 $X=173690 $Y=304400
X725 1 411 130 ICV_7 $T=175260 269280 0 0 $X=175070 $Y=269040
X726 1 133 406 ICV_7 $T=178480 263840 0 0 $X=178290 $Y=263600
X727 1 413 131 ICV_7 $T=178940 280160 0 0 $X=178750 $Y=279920
X728 1 414 406 ICV_7 $T=179860 274720 0 0 $X=179670 $Y=274480
X729 1 125 416 ICV_7 $T=180320 301920 0 0 $X=180130 $Y=301680
X730 1 127 111 ICV_7 $T=181700 296480 1 0 $X=181510 $Y=293520
X731 1 402 137 ICV_7 $T=182160 269280 1 0 $X=181970 $Y=266320
X732 1 412 118 ICV_7 $T=183080 296480 0 0 $X=182890 $Y=296240
X733 1 127 129 ICV_7 $T=184000 301920 0 0 $X=183810 $Y=301680
X734 1 406 418 ICV_7 $T=191820 269280 1 0 $X=191630 $Y=266320
X735 1 402 134 ICV_7 $T=195040 269280 0 0 $X=194850 $Y=269040
X736 1 138 422 ICV_7 $T=195960 301920 0 0 $X=195770 $Y=301680
X737 1 111 118 ICV_7 $T=198260 285600 0 0 $X=198070 $Y=285360
X738 1 142 147 ICV_7 $T=198260 291040 0 0 $X=198070 $Y=290800
X739 1 5 149 ICV_7 $T=203320 263840 0 0 $X=203130 $Y=263600
X740 1 5 427 ICV_7 $T=203320 280160 0 0 $X=203130 $Y=279920
X741 1 151 151 ICV_7 $T=203320 307360 0 0 $X=203130 $Y=307120
X742 1 93 142 ICV_7 $T=205160 301920 0 0 $X=204970 $Y=301680
X743 1 153 141 ICV_7 $T=205620 269280 0 0 $X=205430 $Y=269040
X744 1 425 428 ICV_7 $T=205620 296480 0 0 $X=205430 $Y=296240
X745 1 151 161 ICV_7 $T=213900 291040 0 0 $X=213710 $Y=290800
X746 1 429 7 ICV_7 $T=214360 307360 0 0 $X=214170 $Y=307120
X747 1 434 152 ICV_7 $T=215740 280160 0 0 $X=215550 $Y=279920
X748 1 430 147 ICV_7 $T=217580 291040 1 0 $X=217390 $Y=288080
X749 1 437 159 ICV_7 $T=218040 307360 0 0 $X=217850 $Y=307120
X750 1 436 166 ICV_7 $T=223100 301920 1 0 $X=222910 $Y=298960
X751 1 5 440 ICV_7 $T=224020 274720 0 0 $X=223830 $Y=274480
X752 1 167 439 ICV_7 $T=224940 301920 0 0 $X=224750 $Y=301680
X753 1 5 442 ICV_7 $T=226320 280160 0 0 $X=226130 $Y=279920
X754 1 449 444 ICV_7 $T=245640 285600 1 0 $X=245450 $Y=282640
X755 1 451 180 ICV_7 $T=251620 274720 0 0 $X=251430 $Y=274480
X756 1 179 456 ICV_7 $T=251620 280160 0 0 $X=251430 $Y=279920
X757 1 179 460 ICV_7 $T=254380 269280 0 0 $X=254190 $Y=269040
X758 1 181 122 ICV_7 $T=254380 285600 0 0 $X=254190 $Y=285360
X759 1 458 5 ICV_7 $T=254380 296480 0 0 $X=254190 $Y=296240
X760 1 184 182 ICV_7 $T=255300 301920 1 0 $X=255110 $Y=298960
X761 1 181 457 ICV_7 $T=256680 296480 1 0 $X=256490 $Y=293520
X762 1 462 463 ICV_7 $T=259440 280160 0 0 $X=259250 $Y=279920
X763 1 426 465 ICV_7 $T=261740 291040 0 0 $X=261550 $Y=290800
X764 1 462 186 ICV_7 $T=262200 269280 1 0 $X=262010 $Y=266320
X765 1 172 182 ICV_7 $T=262660 307360 1 0 $X=262470 $Y=304400
X766 1 463 183 ICV_7 $T=265880 285600 0 0 $X=265690 $Y=285360
X767 1 466 190 ICV_7 $T=267260 269280 1 0 $X=267070 $Y=266320
X768 1 467 124 ICV_7 $T=268640 291040 0 0 $X=268450 $Y=290800
X769 1 5 471 ICV_7 $T=274620 285600 0 0 $X=274430 $Y=285360
X770 1 462 186 ICV_7 $T=278760 269280 0 0 $X=278570 $Y=269040
X771 1 197 198 ICV_7 $T=281060 301920 1 0 $X=280870 $Y=298960
X772 1 473 139 ICV_7 $T=282440 269280 0 0 $X=282250 $Y=269040
X773 1 476 426 ICV_7 $T=282440 274720 0 0 $X=282250 $Y=274480
X774 1 426 198 ICV_7 $T=282440 291040 0 0 $X=282250 $Y=290800
X775 1 477 159 ICV_7 $T=282440 307360 0 0 $X=282250 $Y=307120
X776 1 473 190 ICV_7 $T=284740 274720 1 0 $X=284550 $Y=271760
X777 1 202 5 ICV_7 $T=287500 263840 0 0 $X=287310 $Y=263600
X778 1 190 479 ICV_7 $T=290720 280160 0 0 $X=290530 $Y=279920
X779 1 207 483 ICV_7 $T=291180 307360 1 0 $X=290990 $Y=304400
X780 1 472 482 ICV_7 $T=291640 301920 1 0 $X=291450 $Y=298960
X781 1 472 212 ICV_7 $T=296700 307360 1 0 $X=296510 $Y=304400
X782 1 486 211 ICV_7 $T=297160 269280 0 0 $X=296970 $Y=269040
X783 1 209 210 ICV_7 $T=297160 301920 0 0 $X=296970 $Y=301680
X784 1 200 192 ICV_7 $T=300380 280160 0 0 $X=300190 $Y=279920
X785 1 213 218 ICV_7 $T=300840 269280 0 0 $X=300650 $Y=269040
X786 1 488 489 ICV_7 $T=300840 291040 0 0 $X=300650 $Y=290800
X787 1 214 485 ICV_7 $T=300840 296480 0 0 $X=300650 $Y=296240
X788 1 480 216 ICV_7 $T=301760 280160 1 0 $X=301570 $Y=277200
X789 1 217 492 ICV_7 $T=302680 263840 0 0 $X=302490 $Y=263600
X790 1 190 494 ICV_7 $T=304520 269280 1 0 $X=304330 $Y=266320
X791 1 198 204 ICV_7 $T=304520 291040 0 0 $X=304330 $Y=290800
X792 1 222 459 ICV_7 $T=305440 285600 0 0 $X=305250 $Y=285360
X793 1 216 494 ICV_7 $T=307280 274720 0 0 $X=307090 $Y=274480
X794 1 485 223 ICV_7 $T=311880 296480 1 0 $X=311690 $Y=293520
X795 1 497 485 ICV_7 $T=316480 301920 1 0 $X=316290 $Y=298960
X796 1 498 232 ICV_7 $T=320620 307360 0 0 $X=320430 $Y=307120
X797 1 5 3 ICV_7 $T=324300 274720 0 0 $X=324110 $Y=274480
X798 1 5 3 ICV_7 $T=324300 301920 0 0 $X=324110 $Y=301680
X799 1 5 3 ICV_7 $T=324300 307360 0 0 $X=324110 $Y=307120
X800 1 3 5 ICV_7 $T=332120 296480 0 0 $X=331930 $Y=296240
X801 1 3 5 ICV_7 $T=332580 285600 0 0 $X=332390 $Y=285360
X802 1 3 5 ICV_7 $T=333040 291040 0 0 $X=332850 $Y=290800
X803 1 3 5 ICV_7 $T=333500 280160 0 0 $X=333310 $Y=279920
X804 1 3 5 ICV_7 $T=334880 263840 0 0 $X=334690 $Y=263600
X805 1 2 3 4 5 2 11 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 269280 0 0 $X=7630 $Y=269040
X806 1 2 3 317 5 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 274720 0 0 $X=7630 $Y=274480
X807 1 2 3 318 5 2 13 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 280160 0 0 $X=7630 $Y=279920
X808 1 2 3 6 5 2 14 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 301920 0 0 $X=7630 $Y=301680
X809 1 2 3 7 5 2 15 1 sky130_fd_sc_hd__dfrtp_4 $T=8280 307360 0 0 $X=8090 $Y=307120
X810 1 2 3 8 5 2 16 1 sky130_fd_sc_hd__dfrtp_4 $T=9660 285600 0 0 $X=9470 $Y=285360
X811 1 2 3 319 5 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=10120 296480 0 0 $X=9930 $Y=296240
X812 1 2 3 10 5 2 21 1 sky130_fd_sc_hd__dfrtp_4 $T=12880 263840 0 0 $X=12690 $Y=263600
X813 1 2 3 19 5 2 25 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 280160 1 0 $X=20970 $Y=277200
X814 1 2 3 322 5 2 30 1 sky130_fd_sc_hd__dfrtp_4 $T=22540 285600 1 0 $X=22350 $Y=282640
X815 1 2 502 323 5 2 322 1 sky130_fd_sc_hd__dfrtp_4 $T=27140 296480 1 0 $X=26950 $Y=293520
X816 1 2 503 31 5 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 263840 0 0 $X=34770 $Y=263600
X817 1 2 504 325 5 2 22 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 280160 0 0 $X=34770 $Y=279920
X818 1 2 505 327 5 2 39 1 sky130_fd_sc_hd__dfrtp_4 $T=38180 291040 0 0 $X=37990 $Y=290800
X819 1 2 506 345 5 2 60 1 sky130_fd_sc_hd__dfrtp_4 $T=55660 269280 1 0 $X=55470 $Y=266320
X820 1 2 507 349 5 2 319 1 sky130_fd_sc_hd__dfrtp_4 $T=63940 296480 0 0 $X=63750 $Y=296240
X821 1 2 508 355 5 2 320 1 sky130_fd_sc_hd__dfrtp_4 $T=72220 285600 0 0 $X=72030 $Y=285360
X822 1 2 509 356 5 2 65 1 sky130_fd_sc_hd__dfrtp_4 $T=77280 269280 1 0 $X=77090 $Y=266320
X823 1 2 510 367 5 2 74 1 sky130_fd_sc_hd__dfrtp_4 $T=91080 301920 0 0 $X=90890 $Y=301680
X824 1 2 511 375 5 2 317 1 sky130_fd_sc_hd__dfrtp_4 $T=101660 291040 0 0 $X=101470 $Y=290800
X825 1 2 512 96 5 2 100 1 sky130_fd_sc_hd__dfrtp_4 $T=125120 307360 0 0 $X=124930 $Y=307120
X826 1 2 513 387 5 2 103 1 sky130_fd_sc_hd__dfrtp_4 $T=126040 285600 0 0 $X=125850 $Y=285360
X827 1 2 514 388 5 2 102 1 sky130_fd_sc_hd__dfrtp_4 $T=126500 291040 0 0 $X=126310 $Y=290800
X828 1 2 515 391 5 2 99 1 sky130_fd_sc_hd__dfrtp_4 $T=129720 274720 0 0 $X=129530 $Y=274480
X829 1 2 516 400 5 2 123 1 sky130_fd_sc_hd__dfrtp_4 $T=153640 274720 0 0 $X=153450 $Y=274480
X830 1 2 517 404 5 2 128 1 sky130_fd_sc_hd__dfrtp_4 $T=161460 307360 1 0 $X=161270 $Y=304400
X831 1 2 518 407 5 2 321 1 sky130_fd_sc_hd__dfrtp_4 $T=165140 296480 1 0 $X=164950 $Y=293520
X832 1 2 519 417 5 2 140 1 sky130_fd_sc_hd__dfrtp_4 $T=183080 285600 0 0 $X=182890 $Y=285360
X833 1 2 520 419 5 2 146 1 sky130_fd_sc_hd__dfrtp_4 $T=189520 301920 1 0 $X=189330 $Y=298960
X834 1 2 521 427 5 2 145 1 sky130_fd_sc_hd__dfrtp_4 $T=201020 285600 1 0 $X=200830 $Y=282640
X835 1 2 522 149 5 2 153 1 sky130_fd_sc_hd__dfrtp_4 $T=201940 269280 1 0 $X=201750 $Y=266320
X836 1 2 523 440 5 2 168 1 sky130_fd_sc_hd__dfrtp_4 $T=224020 280160 1 0 $X=223830 $Y=277200
X837 1 2 524 441 5 2 171 1 sky130_fd_sc_hd__dfrtp_4 $T=226780 269280 1 0 $X=226590 $Y=266320
X838 1 2 525 443 5 2 446 1 sky130_fd_sc_hd__dfrtp_4 $T=229540 301920 1 0 $X=229350 $Y=298960
X839 1 2 526 447 5 2 177 1 sky130_fd_sc_hd__dfrtp_4 $T=236440 280160 0 0 $X=236250 $Y=279920
X840 1 2 527 176 5 2 178 1 sky130_fd_sc_hd__dfrtp_4 $T=238740 263840 0 0 $X=238550 $Y=263600
X841 1 2 528 449 5 2 183 1 sky130_fd_sc_hd__dfrtp_4 $T=245640 291040 1 0 $X=245450 $Y=288080
X842 1 2 529 454 5 2 185 1 sky130_fd_sc_hd__dfrtp_4 $T=250700 269280 1 0 $X=250510 $Y=266320
X843 1 2 530 457 5 2 465 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 296480 0 0 $X=259250 $Y=296240
X844 1 2 531 466 5 2 193 1 sky130_fd_sc_hd__dfrtp_4 $T=267260 269280 0 0 $X=267070 $Y=269040
X845 1 2 532 191 5 2 468 1 sky130_fd_sc_hd__dfrtp_4 $T=269100 307360 0 0 $X=268910 $Y=307120
X846 1 2 533 471 5 2 318 1 sky130_fd_sc_hd__dfrtp_4 $T=273700 291040 1 0 $X=273510 $Y=288080
X847 1 2 534 481 5 2 215 1 sky130_fd_sc_hd__dfrtp_4 $T=291180 263840 0 0 $X=290990 $Y=263600
X848 1 2 535 492 5 2 229 1 sky130_fd_sc_hd__dfrtp_4 $T=308200 269280 1 0 $X=308010 $Y=266320
X849 1 2 536 496 5 2 231 1 sky130_fd_sc_hd__dfrtp_4 $T=313260 274720 1 0 $X=313070 $Y=271760
X850 1 2 3 234 5 2 239 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 274720 0 0 $X=327790 $Y=274480
X851 1 2 3 235 5 2 240 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 301920 0 0 $X=327790 $Y=301680
X852 1 2 3 233 5 2 241 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 307360 0 0 $X=327790 $Y=307120
X853 1 2 3 446 5 2 247 1 sky130_fd_sc_hd__dfrtp_4 $T=333500 285600 1 0 $X=333310 $Y=282640
X854 1 2 3 237 5 2 248 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 269280 1 0 $X=334690 $Y=266320
X855 1 2 3 238 5 2 249 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 274720 1 0 $X=334690 $Y=271760
X856 1 2 3 318 ICV_8 $T=7820 280160 1 0 $X=7630 $Y=277200
X857 1 2 5 9 ICV_8 $T=10120 291040 1 0 $X=9930 $Y=288080
X858 1 2 5 319 ICV_8 $T=10120 296480 1 0 $X=9930 $Y=293520
X859 1 2 45 45 ICV_8 $T=50600 296480 0 0 $X=50410 $Y=296240
X860 1 2 45 41 ICV_8 $T=51980 301920 1 0 $X=51790 $Y=298960
X861 1 2 344 39 ICV_8 $T=53360 285600 0 0 $X=53170 $Y=285360
X862 1 2 361 368 ICV_8 $T=92000 296480 1 0 $X=91810 $Y=293520
X863 1 2 5 378 ICV_8 $T=106720 285600 0 0 $X=106530 $Y=285360
X864 1 2 384 75 ICV_8 $T=121440 274720 1 0 $X=121250 $Y=271760
X865 1 2 85 101 ICV_8 $T=132480 280160 0 0 $X=132290 $Y=279920
X866 1 2 104 118 ICV_8 $T=149960 307360 1 0 $X=149770 $Y=304400
X867 1 2 399 115 ICV_8 $T=154100 296480 0 0 $X=153910 $Y=296240
X868 1 2 364 401 ICV_8 $T=165140 285600 1 0 $X=164950 $Y=282640
X869 1 2 402 409 ICV_8 $T=169740 269280 1 0 $X=169550 $Y=266320
X870 1 2 5 419 ICV_8 $T=189520 296480 0 0 $X=189330 $Y=296240
X871 1 2 162 445 ICV_8 $T=239660 301920 0 0 $X=239470 $Y=301680
X872 1 2 475 478 ICV_8 $T=287500 291040 0 0 $X=287310 $Y=290800
X873 1 2 481 484 ICV_8 $T=291180 269280 1 0 $X=290990 $Y=266320
X874 1 2 483 459 ICV_8 $T=291640 296480 1 0 $X=291450 $Y=293520
X875 1 2 3 9 17 5 ICV_11 $T=10120 291040 0 0 $X=9930 $Y=290800
X876 1 2 3 320 24 5 ICV_11 $T=21160 274720 1 0 $X=20970 $Y=271760
X877 1 2 3 321 26 5 ICV_11 $T=21160 291040 1 0 $X=20970 $Y=288080
X878 1 2 3 20 27 5 ICV_11 $T=21160 307360 1 0 $X=20970 $Y=304400
X879 1 2 3 22 28 5 ICV_11 $T=22080 269280 1 0 $X=21890 $Y=266320
X880 1 2 537 366 70 5 ICV_11 $T=85100 274720 1 0 $X=84910 $Y=271760
X881 1 2 538 378 90 5 ICV_11 $T=106720 291040 1 0 $X=106530 $Y=288080
X882 1 2 539 394 117 5 ICV_11 $T=143520 291040 1 0 $X=143330 $Y=288080
X883 1 2 540 397 119 5 ICV_11 $T=143980 280160 1 0 $X=143790 $Y=277200
X884 1 2 541 424 150 5 ICV_11 $T=195500 280160 1 0 $X=195310 $Y=277200
X885 1 2 542 442 169 5 ICV_11 $T=225860 285600 1 0 $X=225670 $Y=282640
X886 1 2 543 493 500 5 ICV_11 $T=315560 285600 0 0 $X=315370 $Y=285360
X887 1 2 544 497 501 5 ICV_11 $T=316020 296480 0 0 $X=315830 $Y=296240
X888 1 2 3 465 242 5 ICV_11 $T=332120 280160 1 0 $X=331930 $Y=277200
X889 1 2 3 500 243 5 ICV_11 $T=332120 301920 1 0 $X=331930 $Y=298960
X890 1 2 3 468 244 5 ICV_11 $T=332580 291040 1 0 $X=332390 $Y=288080
X891 1 2 3 501 245 5 ICV_11 $T=333040 296480 1 0 $X=332850 $Y=293520
X892 1 2 3 236 246 5 ICV_11 $T=333040 307360 1 0 $X=332850 $Y=304400
X893 1 2 346 ICV_12 $T=58420 280160 1 0 $X=58230 $Y=277200
X894 1 2 55 ICV_12 $T=65320 274720 0 0 $X=65130 $Y=274480
X895 1 2 363 ICV_12 $T=87400 285600 0 0 $X=87210 $Y=285360
X896 1 2 375 ICV_12 $T=101660 291040 1 0 $X=101470 $Y=288080
X897 1 2 383 ICV_12 $T=119140 296480 0 0 $X=118950 $Y=296240
X898 1 2 391 ICV_12 $T=129720 274720 1 0 $X=129530 $Y=271760
X899 1 2 399 ICV_12 $T=176640 280160 0 0 $X=176450 $Y=279920
X900 1 2 115 ICV_12 $T=177560 274720 0 0 $X=177370 $Y=274480
X901 1 2 420 ICV_12 $T=203320 269280 0 0 $X=203130 $Y=269040
X902 1 2 451 ICV_12 $T=249320 285600 1 0 $X=249130 $Y=282640
X903 1 2 181 ICV_12 $T=253000 307360 1 0 $X=252810 $Y=304400
X904 1 2 200 ICV_12 $T=283820 280160 0 0 $X=283630 $Y=279920
X905 1 2 196 ICV_12 $T=298540 291040 0 0 $X=298350 $Y=290800
X906 1 2 227 ICV_12 $T=322000 301920 0 0 $X=321810 $Y=301680
X907 1 2 234 ICV_12 $T=329820 274720 1 0 $X=329630 $Y=271760
X908 1 2 235 ICV_12 $T=329820 301920 1 0 $X=329630 $Y=298960
X909 1 2 324 ICV_13 $T=31280 301920 1 0 $X=31090 $Y=298960
X910 1 2 32 ICV_13 $T=34040 285600 0 0 $X=33850 $Y=285360
X911 1 2 330 ICV_13 $T=39560 296480 0 0 $X=39370 $Y=296240
X912 1 2 334 ICV_13 $T=44160 269280 1 0 $X=43970 $Y=266320
X913 1 2 44 ICV_13 $T=48760 291040 0 0 $X=48570 $Y=290800
X914 1 2 46 ICV_13 $T=48760 307360 0 0 $X=48570 $Y=307120
X915 1 2 29 ICV_13 $T=57960 307360 0 0 $X=57770 $Y=307120
X916 1 2 5 ICV_13 $T=68540 285600 0 0 $X=68350 $Y=285360
X917 1 2 355 ICV_13 $T=70380 285600 1 0 $X=70190 $Y=282640
X918 1 2 368 ICV_13 $T=84640 301920 1 0 $X=84450 $Y=298960
X919 1 2 43 ICV_13 $T=86020 296480 0 0 $X=85830 $Y=296240
X920 1 2 67 ICV_13 $T=90160 307360 0 0 $X=89970 $Y=307120
X921 1 2 98 ICV_13 $T=127880 269280 0 0 $X=127690 $Y=269040
X922 1 2 361 ICV_13 $T=128340 296480 1 0 $X=128150 $Y=293520
X923 1 2 351 ICV_13 $T=146280 280160 0 0 $X=146090 $Y=279920
X924 1 2 124 ICV_13 $T=162380 296480 0 0 $X=162190 $Y=296240
X925 1 2 410 ICV_13 $T=170200 296480 0 0 $X=170010 $Y=296240
X926 1 2 129 ICV_13 $T=170200 307360 0 0 $X=170010 $Y=307120
X927 1 2 129 ICV_13 $T=171120 301920 1 0 $X=170930 $Y=298960
X928 1 2 93 ICV_13 $T=182160 307360 0 0 $X=181970 $Y=307120
X929 1 2 424 ICV_13 $T=189980 274720 0 0 $X=189790 $Y=274480
X930 1 2 431 ICV_13 $T=203320 291040 1 0 $X=203130 $Y=288080
X931 1 2 156 ICV_13 $T=208380 263840 0 0 $X=208190 $Y=263600
X932 1 2 431 ICV_13 $T=211140 285600 0 0 $X=210950 $Y=285360
X933 1 2 142 ICV_13 $T=216660 301920 1 0 $X=216470 $Y=298960
X934 1 2 439 ICV_13 $T=216660 307360 1 0 $X=216470 $Y=304400
X935 1 2 163 ICV_13 $T=217580 263840 0 0 $X=217390 $Y=263600
X936 1 2 443 ICV_13 $T=227700 296480 1 0 $X=227510 $Y=293520
X937 1 2 43 ICV_13 $T=254380 301920 0 0 $X=254190 $Y=301680
X938 1 2 188 ICV_13 $T=258520 274720 1 0 $X=258330 $Y=271760
X939 1 2 5 ICV_13 $T=263580 269280 0 0 $X=263390 $Y=269040
X940 1 2 444 ICV_13 $T=268640 285600 0 0 $X=268450 $Y=285360
X941 1 2 472 ICV_13 $T=276460 291040 0 0 $X=276270 $Y=290800
X942 1 2 201 ICV_13 $T=282440 285600 0 0 $X=282250 $Y=285360
X943 1 2 210 ICV_13 $T=296700 274720 1 0 $X=296510 $Y=271760
X944 1 2 216 ICV_13 $T=299920 307360 0 0 $X=299730 $Y=307120
X945 1 2 490 ICV_13 $T=300840 296480 1 0 $X=300650 $Y=293520
X946 1 2 216 ICV_13 $T=308200 307360 1 0 $X=308010 $Y=304400
X947 1 2 210 ICV_13 $T=310040 307360 0 0 $X=309850 $Y=307120
X948 1 2 226 ICV_13 $T=310500 301920 0 0 $X=310310 $Y=301680
X949 1 2 ICV_14 $T=19780 269280 1 0 $X=19590 $Y=266320
X950 1 2 ICV_14 $T=19780 285600 1 0 $X=19590 $Y=282640
X951 1 2 ICV_14 $T=33580 291040 0 0 $X=33390 $Y=290800
X952 1 2 ICV_14 $T=47840 269280 1 0 $X=47650 $Y=266320
X953 1 2 ICV_14 $T=47840 280160 1 0 $X=47650 $Y=277200
X954 1 2 ICV_14 $T=47840 285600 1 0 $X=47650 $Y=282640
X955 1 2 ICV_14 $T=47840 296480 1 0 $X=47650 $Y=293520
X956 1 2 ICV_14 $T=61640 296480 0 0 $X=61450 $Y=296240
X957 1 2 ICV_14 $T=75900 301920 1 0 $X=75710 $Y=298960
X958 1 2 ICV_14 $T=89700 285600 0 0 $X=89510 $Y=285360
X959 1 2 ICV_14 $T=103960 280160 1 0 $X=103770 $Y=277200
X960 1 2 ICV_14 $T=103960 291040 1 0 $X=103770 $Y=288080
X961 1 2 ICV_14 $T=117760 274720 0 0 $X=117570 $Y=274480
X962 1 2 ICV_14 $T=117760 301920 0 0 $X=117570 $Y=301680
X963 1 2 ICV_14 $T=132020 307360 1 0 $X=131830 $Y=304400
X964 1 2 ICV_14 $T=145820 301920 0 0 $X=145630 $Y=301680
X965 1 2 ICV_14 $T=145820 307360 0 0 $X=145630 $Y=307120
X966 1 2 ICV_14 $T=160080 285600 1 0 $X=159890 $Y=282640
X967 1 2 ICV_14 $T=173880 280160 0 0 $X=173690 $Y=279920
X968 1 2 ICV_14 $T=173880 296480 0 0 $X=173690 $Y=296240
X969 1 2 ICV_14 $T=230000 269280 0 0 $X=229810 $Y=269040
X970 1 2 ICV_14 $T=272320 269280 1 0 $X=272130 $Y=266320
X971 1 2 ICV_14 $T=272320 280160 1 0 $X=272130 $Y=277200
X972 1 2 ICV_14 $T=286120 274720 0 0 $X=285930 $Y=274480
X973 1 5 ICV_15 $T=31740 263840 0 0 $X=31550 $Y=263600
X974 1 5 ICV_15 $T=31740 280160 0 0 $X=31550 $Y=279920
X975 1 29 ICV_15 $T=31740 296480 0 0 $X=31550 $Y=296240
X976 1 339 ICV_15 $T=46000 274720 1 0 $X=45810 $Y=271760
X977 1 328 ICV_15 $T=46000 291040 1 0 $X=45810 $Y=288080
X978 1 52 ICV_15 $T=59800 274720 0 0 $X=59610 $Y=274480
X979 1 53 ICV_15 $T=59800 301920 0 0 $X=59610 $Y=301680
X980 1 90 ICV_15 $T=115920 285600 0 0 $X=115730 $Y=285360
X981 1 79 ICV_15 $T=115920 291040 0 0 $X=115730 $Y=290800
X982 1 392 ICV_15 $T=130180 291040 1 0 $X=129990 $Y=288080
X983 1 109 ICV_15 $T=143980 263840 0 0 $X=143790 $Y=263600
X984 1 5 ICV_15 $T=143980 274720 0 0 $X=143790 $Y=274480
X985 1 402 ICV_15 $T=158240 274720 1 0 $X=158050 $Y=271760
X986 1 321 ICV_15 $T=172040 291040 0 0 $X=171850 $Y=290800
X987 1 421 ICV_15 $T=186300 274720 1 0 $X=186110 $Y=271760
X988 1 422 ICV_15 $T=186300 301920 1 0 $X=186110 $Y=298960
X989 1 426 ICV_15 $T=200100 296480 0 0 $X=199910 $Y=296240
X990 1 147 ICV_15 $T=214360 285600 1 0 $X=214170 $Y=282640
X991 1 433 ICV_15 $T=214360 291040 1 0 $X=214170 $Y=288080
X992 1 142 ICV_15 $T=214360 296480 1 0 $X=214170 $Y=293520
X993 1 5 ICV_15 $T=228160 296480 0 0 $X=227970 $Y=296240
X994 1 211 ICV_15 $T=298540 280160 1 0 $X=298350 $Y=277200
X995 1 487 ICV_15 $T=298540 301920 1 0 $X=298350 $Y=298960
X996 1 5 ICV_15 $T=312340 269280 0 0 $X=312150 $Y=269040
X997 1 5 ICV_15 $T=312340 285600 0 0 $X=312150 $Y=285360
X998 1 233 ICV_15 $T=326600 307360 1 0 $X=326410 $Y=304400
X999 1 2 317 ICV_16 $T=11500 274720 1 0 $X=11310 $Y=271760
X1000 1 2 8 ICV_16 $T=11500 285600 1 0 $X=11310 $Y=282640
X1001 1 2 6 ICV_16 $T=11500 301920 1 0 $X=11310 $Y=298960
X1002 1 2 7 ICV_16 $T=11960 307360 1 0 $X=11770 $Y=304400
X1003 1 2 10 ICV_16 $T=12880 269280 1 0 $X=12690 $Y=266320
X1004 1 2 19 ICV_16 $T=23920 274720 0 0 $X=23730 $Y=274480
X1005 1 2 23 ICV_16 $T=23920 307360 0 0 $X=23730 $Y=307120
X1006 1 2 320 ICV_16 $T=24380 269280 0 0 $X=24190 $Y=269040
X1007 1 2 321 ICV_16 $T=24840 285600 0 0 $X=24650 $Y=285360
X1008 1 2 20 ICV_16 $T=24840 301920 0 0 $X=24650 $Y=301680
X1009 1 2 329 ICV_16 $T=39100 274720 1 0 $X=38910 $Y=271760
X1010 1 2 331 ICV_16 $T=56580 291040 1 0 $X=56390 $Y=288080
X1011 1 2 349 ICV_16 $T=63940 301920 1 0 $X=63750 $Y=298960
X1012 1 2 45 ICV_16 $T=68080 307360 1 0 $X=67890 $Y=304400
X1013 1 2 362 ICV_16 $T=79580 301920 0 0 $X=79390 $Y=301680
X1014 1 2 62 ICV_16 $T=80040 274720 0 0 $X=79850 $Y=274480
X1015 1 2 320 ICV_16 $T=80040 280160 0 0 $X=79850 $Y=279920
X1016 1 2 365 ICV_16 $T=85100 285600 1 0 $X=84910 $Y=282640
X1017 1 2 69 ICV_16 $T=94760 301920 1 0 $X=94570 $Y=298960
X1018 1 2 70 ICV_16 $T=95680 280160 1 0 $X=95490 $Y=277200
X1019 1 2 380 ICV_16 $T=109940 280160 0 0 $X=109750 $Y=279920
X1020 1 2 88 ICV_16 $T=120520 301920 0 0 $X=120330 $Y=301680
X1021 1 2 386 ICV_16 $T=133400 269280 1 0 $X=133210 $Y=266320
X1022 1 2 99 ICV_16 $T=133400 274720 1 0 $X=133210 $Y=271760
X1023 1 2 100 ICV_16 $T=134320 301920 0 0 $X=134130 $Y=301680
X1024 1 2 120 ICV_16 $T=161460 263840 0 0 $X=161270 $Y=263600
X1025 1 2 399 ICV_16 $T=180320 291040 0 0 $X=180130 $Y=290800
X1026 1 2 140 ICV_16 $T=189060 280160 0 0 $X=188870 $Y=279920
X1027 1 2 141 ICV_16 $T=195040 263840 0 0 $X=194850 $Y=263600
X1028 1 2 432 ICV_16 $T=207000 280160 0 0 $X=206810 $Y=279920
X1029 1 2 155 ICV_16 $T=208840 301920 0 0 $X=208650 $Y=301680
X1030 1 2 433 ICV_16 $T=221260 291040 1 0 $X=221070 $Y=288080
X1031 1 2 445 ICV_16 $T=231380 291040 0 0 $X=231190 $Y=290800
X1032 1 2 171 ICV_16 $T=232760 274720 1 0 $X=232570 $Y=271760
X1033 1 2 446 ICV_16 $T=233680 296480 1 0 $X=233490 $Y=293520
X1034 1 2 447 ICV_16 $T=236440 280160 1 0 $X=236250 $Y=277200
X1035 1 2 177 ICV_16 $T=244720 274720 0 0 $X=244530 $Y=274480
X1036 1 2 450 ICV_16 $T=246100 291040 0 0 $X=245910 $Y=290800
X1037 1 2 186 ICV_16 $T=259900 280160 1 0 $X=259710 $Y=277200
X1038 1 2 461 ICV_16 $T=263120 280160 0 0 $X=262930 $Y=279920
X1039 1 2 470 ICV_16 $T=274620 280160 1 0 $X=274430 $Y=277200
X1040 1 2 495 ICV_16 $T=306820 285600 1 0 $X=306630 $Y=282640
X1041 1 2 493 ICV_16 $T=314640 291040 1 0 $X=314450 $Y=288080
X1042 1 2 501 ICV_16 $T=318780 291040 0 0 $X=318590 $Y=290800
X1043 1 2 227 ICV_16 $T=319240 307360 1 0 $X=319050 $Y=304400
X1044 1 2 231 ICV_16 $T=319700 269280 1 0 $X=319510 $Y=266320
X1045 1 2 499 ICV_16 $T=320160 301920 1 0 $X=319970 $Y=298960
X1046 1 2 496 ICV_16 $T=321540 269280 0 0 $X=321350 $Y=269040
X1047 1 2 500 ICV_16 $T=335800 296480 0 0 $X=335610 $Y=296240
X1048 1 2 322 2 328 1 sky130_fd_sc_hd__inv_8 $T=35420 296480 0 0 $X=35230 $Y=296240
X1049 1 2 22 2 331 1 sky130_fd_sc_hd__inv_8 $T=37720 285600 0 0 $X=37530 $Y=285360
X1050 1 2 36 2 334 1 sky130_fd_sc_hd__inv_8 $T=40020 269280 1 0 $X=39830 $Y=266320
X1051 1 2 39 2 343 1 sky130_fd_sc_hd__inv_8 $T=48300 285600 0 0 $X=48110 $Y=285360
X1052 1 2 319 2 357 1 sky130_fd_sc_hd__inv_8 $T=71760 301920 0 0 $X=71570 $Y=301680
X1053 1 2 65 2 350 1 sky130_fd_sc_hd__inv_8 $T=78200 263840 0 0 $X=78010 $Y=263600
X1054 1 2 320 2 363 1 sky130_fd_sc_hd__inv_8 $T=80040 285600 1 0 $X=79850 $Y=282640
X1055 1 2 69 2 368 1 sky130_fd_sc_hd__inv_8 $T=90620 307360 1 0 $X=90430 $Y=304400
X1056 1 2 70 2 372 1 sky130_fd_sc_hd__inv_8 $T=94300 274720 0 0 $X=94110 $Y=274480
X1057 1 2 9 2 72 1 sky130_fd_sc_hd__inv_8 $T=94760 263840 0 0 $X=94570 $Y=263600
X1058 1 2 74 2 86 1 sky130_fd_sc_hd__inv_8 $T=104420 301920 0 0 $X=104230 $Y=301680
X1059 1 2 317 2 381 1 sky130_fd_sc_hd__inv_8 $T=108100 296480 1 0 $X=107910 $Y=293520
X1060 1 2 90 2 382 1 sky130_fd_sc_hd__inv_8 $T=119140 285600 0 0 $X=118950 $Y=285360
X1061 1 2 99 2 384 1 sky130_fd_sc_hd__inv_8 $T=133400 280160 1 0 $X=133210 $Y=277200
X1062 1 2 102 2 390 1 sky130_fd_sc_hd__inv_8 $T=134320 291040 1 0 $X=134130 $Y=288080
X1063 1 2 100 2 104 1 sky130_fd_sc_hd__inv_8 $T=134320 307360 1 0 $X=134130 $Y=304400
X1064 1 2 103 2 110 1 sky130_fd_sc_hd__inv_8 $T=140300 274720 1 0 $X=140110 $Y=271760
X1065 1 2 109 2 113 1 sky130_fd_sc_hd__inv_8 $T=147200 263840 0 0 $X=147010 $Y=263600
X1066 1 2 117 2 396 1 sky130_fd_sc_hd__inv_8 $T=149960 285600 0 0 $X=149770 $Y=285360
X1067 1 2 119 2 401 1 sky130_fd_sc_hd__inv_8 $T=155020 269280 0 0 $X=154830 $Y=269040
X1068 1 2 123 2 409 1 sky130_fd_sc_hd__inv_8 $T=166060 269280 0 0 $X=165870 $Y=269040
X1069 1 2 321 2 410 1 sky130_fd_sc_hd__inv_8 $T=175260 291040 0 0 $X=175070 $Y=290800
X1070 1 2 128 2 132 1 sky130_fd_sc_hd__inv_8 $T=175260 301920 0 0 $X=175070 $Y=301680
X1071 1 2 140 2 418 1 sky130_fd_sc_hd__inv_8 $T=189520 285600 1 0 $X=189330 $Y=282640
X1072 1 2 145 2 425 1 sky130_fd_sc_hd__inv_8 $T=199180 291040 1 0 $X=198990 $Y=288080
X1073 1 2 150 2 420 1 sky130_fd_sc_hd__inv_8 $T=203320 274720 0 0 $X=203130 $Y=274480
X1074 1 2 146 2 422 1 sky130_fd_sc_hd__inv_8 $T=203780 301920 1 0 $X=203590 $Y=298960
X1075 1 2 153 2 158 1 sky130_fd_sc_hd__inv_8 $T=209300 269280 0 0 $X=209110 $Y=269040
X1076 1 2 168 2 431 1 sky130_fd_sc_hd__inv_8 $T=225860 274720 1 0 $X=225670 $Y=271760
X1077 1 2 169 2 433 1 sky130_fd_sc_hd__inv_8 $T=231380 285600 0 0 $X=231190 $Y=285360
X1078 1 2 171 2 174 1 sky130_fd_sc_hd__inv_8 $T=232760 269280 0 0 $X=232570 $Y=269040
X1079 1 2 446 2 439 1 sky130_fd_sc_hd__inv_8 $T=232760 296480 0 0 $X=232570 $Y=296240
X1080 1 2 177 2 451 1 sky130_fd_sc_hd__inv_8 $T=245640 280160 1 0 $X=245450 $Y=277200
X1081 1 2 185 2 188 1 sky130_fd_sc_hd__inv_8 $T=259440 269280 0 0 $X=259250 $Y=269040
X1082 1 2 183 2 463 1 sky130_fd_sc_hd__inv_8 $T=259900 291040 1 0 $X=259710 $Y=288080
X1083 1 2 465 2 452 1 sky130_fd_sc_hd__inv_8 $T=263580 296480 1 0 $X=263390 $Y=293520
X1084 1 2 468 2 458 1 sky130_fd_sc_hd__inv_8 $T=273700 307360 1 0 $X=273510 $Y=304400
X1085 1 2 193 2 473 1 sky130_fd_sc_hd__inv_8 $T=277380 263840 0 0 $X=277190 $Y=263600
X1086 1 2 318 2 475 1 sky130_fd_sc_hd__inv_8 $T=278300 285600 0 0 $X=278110 $Y=285360
X1087 1 2 208 2 483 1 sky130_fd_sc_hd__inv_8 $T=295780 307360 0 0 $X=295590 $Y=307120
X1088 1 2 229 2 228 1 sky130_fd_sc_hd__inv_8 $T=315560 263840 0 0 $X=315370 $Y=263600
X1089 1 2 500 2 479 1 sky130_fd_sc_hd__inv_8 $T=316020 285600 1 0 $X=315830 $Y=282640
X1090 1 2 231 2 494 1 sky130_fd_sc_hd__inv_8 $T=316480 269280 0 0 $X=316290 $Y=269040
X1091 1 2 501 2 489 1 sky130_fd_sc_hd__inv_8 $T=318780 296480 1 0 $X=318590 $Y=293520
X1092 1 2 29 324 2 323 1 sky130_fd_sc_hd__nor2_4 $T=34960 301920 1 0 $X=34770 $Y=298960
X1093 1 2 32 326 2 325 1 sky130_fd_sc_hd__nor2_4 $T=37260 291040 1 0 $X=37070 $Y=288080
X1094 1 2 32 329 2 31 1 sky130_fd_sc_hd__nor2_4 $T=39100 269280 0 0 $X=38910 $Y=269040
X1095 1 2 29 332 2 35 1 sky130_fd_sc_hd__nor2_4 $T=39100 307360 1 0 $X=38910 $Y=304400
X1096 1 2 32 333 2 327 1 sky130_fd_sc_hd__nor2_4 $T=40020 285600 1 0 $X=39830 $Y=282640
X1097 1 2 32 342 2 345 1 sky130_fd_sc_hd__nor2_4 $T=51520 263840 0 0 $X=51330 $Y=263600
X1098 1 2 351 353 2 349 1 sky130_fd_sc_hd__nor2_4 $T=68080 296480 1 0 $X=67890 $Y=293520
X1099 1 2 64 352 2 356 1 sky130_fd_sc_hd__nor2_4 $T=77280 274720 1 0 $X=77090 $Y=271760
X1100 1 2 351 358 2 355 1 sky130_fd_sc_hd__nor2_4 $T=77280 291040 0 0 $X=77090 $Y=290800
X1101 1 2 351 360 2 66 1 sky130_fd_sc_hd__nor2_4 $T=80500 301920 1 0 $X=80310 $Y=298960
X1102 1 2 64 369 2 366 1 sky130_fd_sc_hd__nor2_4 $T=90620 280160 1 0 $X=90430 $Y=277200
X1103 1 2 64 371 2 68 1 sky130_fd_sc_hd__nor2_4 $T=92920 269280 1 0 $X=92730 $Y=266320
X1104 1 2 67 71 2 367 1 sky130_fd_sc_hd__nor2_4 $T=93840 307360 0 0 $X=93650 $Y=307120
X1105 1 2 64 373 2 378 1 sky130_fd_sc_hd__nor2_4 $T=103960 280160 0 0 $X=103770 $Y=279920
X1106 1 2 85 379 2 375 1 sky130_fd_sc_hd__nor2_4 $T=108560 296480 0 0 $X=108370 $Y=296240
X1107 1 2 95 389 2 388 1 sky130_fd_sc_hd__nor2_4 $T=124200 296480 1 0 $X=124010 $Y=293520
X1108 1 2 98 386 2 391 1 sky130_fd_sc_hd__nor2_4 $T=131560 269280 0 0 $X=131370 $Y=269040
X1109 1 2 85 101 2 387 1 sky130_fd_sc_hd__nor2_4 $T=133400 285600 1 0 $X=133210 $Y=282640
X1110 1 2 95 392 2 394 1 sky130_fd_sc_hd__nor2_4 $T=133860 296480 1 0 $X=133670 $Y=293520
X1111 1 2 351 398 2 397 1 sky130_fd_sc_hd__nor2_4 $T=149960 280160 0 0 $X=149770 $Y=279920
X1112 1 2 351 405 2 400 1 sky130_fd_sc_hd__nor2_4 $T=161460 274720 1 0 $X=161270 $Y=271760
X1113 1 2 124 408 2 407 1 sky130_fd_sc_hd__nor2_4 $T=166060 296480 0 0 $X=165870 $Y=296240
X1114 1 2 125 126 2 404 1 sky130_fd_sc_hd__nor2_4 $T=166060 307360 0 0 $X=165870 $Y=307120
X1115 1 2 125 415 2 419 1 sky130_fd_sc_hd__nor2_4 $T=180320 307360 1 0 $X=180130 $Y=304400
X1116 1 2 131 413 2 417 1 sky130_fd_sc_hd__nor2_4 $T=182620 280160 0 0 $X=182430 $Y=279920
X1117 1 2 131 423 2 424 1 sky130_fd_sc_hd__nor2_4 $T=193660 274720 0 0 $X=193470 $Y=274480
X1118 1 2 152 432 2 427 1 sky130_fd_sc_hd__nor2_4 $T=207000 291040 1 0 $X=206810 $Y=288080
X1119 1 2 152 434 2 440 1 sky130_fd_sc_hd__nor2_4 $T=218040 285600 1 0 $X=217850 $Y=282640
X1120 1 2 163 164 2 441 1 sky130_fd_sc_hd__nor2_4 $T=221260 263840 0 0 $X=221070 $Y=263600
X1121 1 2 152 438 2 442 1 sky130_fd_sc_hd__nor2_4 $T=221260 280160 0 0 $X=221070 $Y=279920
X1122 1 2 165 437 2 443 1 sky130_fd_sc_hd__nor2_4 $T=222180 307360 0 0 $X=221990 $Y=307120
X1123 1 2 124 448 2 447 1 sky130_fd_sc_hd__nor2_4 $T=240120 291040 0 0 $X=239930 $Y=290800
X1124 1 2 172 453 2 457 1 sky130_fd_sc_hd__nor2_4 $T=250240 307360 0 0 $X=250050 $Y=307120
X1125 1 2 179 456 2 449 1 sky130_fd_sc_hd__nor2_4 $T=251620 285600 1 0 $X=251430 $Y=282640
X1126 1 2 179 460 2 454 1 sky130_fd_sc_hd__nor2_4 $T=254380 274720 1 0 $X=254190 $Y=271760
X1127 1 2 124 467 2 471 1 sky130_fd_sc_hd__nor2_4 $T=272320 291040 0 0 $X=272130 $Y=290800
X1128 1 2 192 470 2 466 1 sky130_fd_sc_hd__nor2_4 $T=274620 274720 0 0 $X=274430 $Y=274480
X1129 1 2 179 194 2 195 1 sky130_fd_sc_hd__nor2_4 $T=275080 269280 1 0 $X=274890 $Y=266320
X1130 1 2 204 477 2 205 1 sky130_fd_sc_hd__nor2_4 $T=287960 307360 0 0 $X=287770 $Y=307120
X1131 1 2 192 484 2 481 1 sky130_fd_sc_hd__nor2_4 $T=292560 274720 1 0 $X=292370 $Y=271760
X1132 1 2 192 480 2 493 1 sky130_fd_sc_hd__nor2_4 $T=301760 285600 1 0 $X=301570 $Y=282640
X1133 1 2 131 217 2 492 1 sky130_fd_sc_hd__nor2_4 $T=306360 263840 0 0 $X=306170 $Y=263600
X1134 1 2 192 495 2 496 1 sky130_fd_sc_hd__nor2_4 $T=306360 280160 0 0 $X=306170 $Y=279920
X1135 1 2 204 490 2 497 1 sky130_fd_sc_hd__nor2_4 $T=306360 296480 0 0 $X=306170 $Y=296240
X1136 1 2 204 498 2 230 1 sky130_fd_sc_hd__nor2_4 $T=315560 307360 0 0 $X=315370 $Y=307120
X1137 1 2 34 37 330 335 2 33 1 sky130_fd_sc_hd__o22a_4 $T=42320 307360 0 0 $X=42130 $Y=307120
X1138 1 2 328 37 330 338 2 324 1 sky130_fd_sc_hd__o22a_4 $T=43240 296480 0 0 $X=43050 $Y=296240
X1139 1 2 334 336 340 339 2 329 1 sky130_fd_sc_hd__o22a_4 $T=49220 274720 1 0 $X=49030 $Y=271760
X1140 1 2 331 37 330 344 2 326 1 sky130_fd_sc_hd__o22a_4 $T=49220 291040 1 0 $X=49030 $Y=288080
X1141 1 2 41 37 330 337 2 332 1 sky130_fd_sc_hd__o22a_4 $T=49220 307360 1 0 $X=49030 $Y=304400
X1142 1 2 343 336 340 341 2 333 1 sky130_fd_sc_hd__o22a_4 $T=50600 280160 0 0 $X=50410 $Y=279920
X1143 1 2 49 336 340 346 2 342 1 sky130_fd_sc_hd__o22a_4 $T=58420 274720 1 0 $X=58230 $Y=271760
X1144 1 2 53 37 330 347 2 51 1 sky130_fd_sc_hd__o22a_4 $T=60720 307360 1 0 $X=60530 $Y=304400
X1145 1 2 61 336 340 348 2 54 1 sky130_fd_sc_hd__o22a_4 $T=63020 269280 0 0 $X=62830 $Y=269040
X1146 1 2 350 336 340 354 2 352 1 sky130_fd_sc_hd__o22a_4 $T=67620 274720 0 0 $X=67430 $Y=274480
X1147 1 2 357 361 359 362 2 353 1 sky130_fd_sc_hd__o22a_4 $T=79580 296480 0 0 $X=79390 $Y=296240
X1148 1 2 363 361 359 365 2 358 1 sky130_fd_sc_hd__o22a_4 $T=82340 291040 1 0 $X=82150 $Y=288080
X1149 1 2 368 361 359 370 2 360 1 sky130_fd_sc_hd__o22a_4 $T=91080 296480 0 0 $X=90890 $Y=296240
X1150 1 2 73 75 377 83 2 371 1 sky130_fd_sc_hd__o22a_4 $T=105340 269280 1 0 $X=105150 $Y=266320
X1151 1 2 372 75 377 376 2 369 1 sky130_fd_sc_hd__o22a_4 $T=105340 274720 1 0 $X=105150 $Y=271760
X1152 1 2 86 82 78 374 2 71 1 sky130_fd_sc_hd__o22a_4 $T=105800 307360 0 0 $X=105610 $Y=307120
X1153 1 2 382 75 377 380 2 373 1 sky130_fd_sc_hd__o22a_4 $T=109940 280160 1 0 $X=109750 $Y=277200
X1154 1 2 381 82 78 383 2 379 1 sky130_fd_sc_hd__o22a_4 $T=111320 301920 1 0 $X=111130 $Y=298960
X1155 1 2 91 75 377 92 2 89 1 sky130_fd_sc_hd__o22a_4 $T=114540 269280 1 0 $X=114350 $Y=266320
X1156 1 2 384 75 377 385 2 386 1 sky130_fd_sc_hd__o22a_4 $T=121440 269280 0 0 $X=121250 $Y=269040
X1157 1 2 390 361 359 393 2 389 1 sky130_fd_sc_hd__o22a_4 $T=132020 296480 0 0 $X=131830 $Y=296240
X1158 1 2 396 361 359 395 2 392 1 sky130_fd_sc_hd__o22a_4 $T=141680 296480 1 0 $X=141490 $Y=293520
X1159 1 2 401 402 406 403 2 398 1 sky130_fd_sc_hd__o22a_4 $T=161920 280160 1 0 $X=161730 $Y=277200
X1160 1 2 409 402 406 411 2 405 1 sky130_fd_sc_hd__o22a_4 $T=169740 274720 1 0 $X=169550 $Y=271760
X1161 1 2 410 127 412 129 2 408 1 sky130_fd_sc_hd__o22a_4 $T=174800 301920 1 0 $X=174610 $Y=298960
X1162 1 2 132 127 129 135 2 126 1 sky130_fd_sc_hd__o22a_4 $T=175720 307360 0 0 $X=175530 $Y=307120
X1163 1 2 133 402 406 137 2 136 1 sky130_fd_sc_hd__o22a_4 $T=182160 263840 0 0 $X=181970 $Y=263600
X1164 1 2 418 402 406 414 2 413 1 sky130_fd_sc_hd__o22a_4 $T=183540 274720 0 0 $X=183350 $Y=274480
X1165 1 2 420 402 406 421 2 423 1 sky130_fd_sc_hd__o22a_4 $T=189520 274720 1 0 $X=189330 $Y=271760
X1166 1 2 422 127 129 416 2 415 1 sky130_fd_sc_hd__o22a_4 $T=189520 307360 1 0 $X=189330 $Y=304400
X1167 1 2 425 147 151 428 2 432 1 sky130_fd_sc_hd__o22a_4 $T=205160 291040 0 0 $X=204970 $Y=290800
X1168 1 2 155 147 151 429 2 154 1 sky130_fd_sc_hd__o22a_4 $T=207000 307360 0 0 $X=206810 $Y=307120
X1169 1 2 431 147 430 151 2 434 1 sky130_fd_sc_hd__o22a_4 $T=214820 285600 0 0 $X=214630 $Y=285360
X1170 1 2 433 147 151 435 2 438 1 sky130_fd_sc_hd__o22a_4 $T=217580 291040 0 0 $X=217390 $Y=290800
X1171 1 2 439 166 167 436 2 437 1 sky130_fd_sc_hd__o22a_4 $T=223100 307360 1 0 $X=222910 $Y=304400
X1172 1 2 451 444 445 450 2 448 1 sky130_fd_sc_hd__o22a_4 $T=246100 285600 0 0 $X=245910 $Y=285360
X1173 1 2 452 182 184 455 2 453 1 sky130_fd_sc_hd__o22a_4 $T=255300 307360 1 0 $X=255110 $Y=304400
X1174 1 2 463 186 462 461 2 456 1 sky130_fd_sc_hd__o22a_4 $T=259440 285600 1 0 $X=259250 $Y=282640
X1175 1 2 458 182 184 187 2 189 1 sky130_fd_sc_hd__o22a_4 $T=259440 307360 0 0 $X=259250 $Y=307120
X1176 1 2 188 186 462 464 2 460 1 sky130_fd_sc_hd__o22a_4 $T=262200 274720 1 0 $X=262010 $Y=271760
X1177 1 2 473 186 462 469 2 470 1 sky130_fd_sc_hd__o22a_4 $T=275540 274720 1 0 $X=275350 $Y=271760
X1178 1 2 475 472 198 478 2 467 1 sky130_fd_sc_hd__o22a_4 $T=281980 296480 1 0 $X=281790 $Y=293520
X1179 1 2 202 186 462 203 2 194 1 sky130_fd_sc_hd__o22a_4 $T=282900 269280 1 0 $X=282710 $Y=266320
X1180 1 2 197 472 198 474 2 199 1 sky130_fd_sc_hd__o22a_4 $T=282900 307360 1 0 $X=282710 $Y=304400
X1181 1 2 479 186 462 476 2 480 1 sky130_fd_sc_hd__o22a_4 $T=289800 280160 1 0 $X=289610 $Y=277200
X1182 1 2 483 472 198 482 2 477 1 sky130_fd_sc_hd__o22a_4 $T=289800 301920 0 0 $X=289610 $Y=301680
X1183 1 2 211 210 216 486 2 484 1 sky130_fd_sc_hd__o22a_4 $T=299920 274720 0 0 $X=299730 $Y=274480
X1184 1 2 209 210 216 487 2 207 1 sky130_fd_sc_hd__o22a_4 $T=301760 307360 1 0 $X=301570 $Y=304400
X1185 1 2 223 472 198 224 2 221 1 sky130_fd_sc_hd__o22a_4 $T=303600 307360 0 0 $X=303410 $Y=307120
X1186 1 2 489 472 198 488 2 490 1 sky130_fd_sc_hd__o22a_4 $T=304520 296480 1 0 $X=304330 $Y=293520
X1187 1 2 494 210 216 491 2 495 1 sky130_fd_sc_hd__o22a_4 $T=306360 280160 1 0 $X=306170 $Y=277200
X1188 1 2 227 210 216 499 2 498 1 sky130_fd_sc_hd__o22a_4 $T=311880 307360 1 0 $X=311690 $Y=304400
X1189 1 2 42 2 32 1 sky130_fd_sc_hd__buf_1 $T=50600 269280 1 0 $X=50410 $Y=266320
X1190 1 2 55 2 336 1 sky130_fd_sc_hd__buf_1 $T=63020 274720 0 0 $X=62830 $Y=274480
X1191 1 2 55 2 37 1 sky130_fd_sc_hd__buf_1 $T=63480 285600 0 0 $X=63290 $Y=285360
X1192 1 2 57 2 330 1 sky130_fd_sc_hd__buf_1 $T=65320 291040 1 0 $X=65130 $Y=288080
X1193 1 2 62 2 45 1 sky130_fd_sc_hd__buf_1 $T=69000 285600 1 0 $X=68810 $Y=282640
X1194 1 2 57 2 340 1 sky130_fd_sc_hd__buf_1 $T=69920 280160 1 0 $X=69730 $Y=277200
X1195 1 2 62 2 47 1 sky130_fd_sc_hd__buf_1 $T=77740 274720 0 0 $X=77550 $Y=274480
X1196 1 2 42 2 64 1 sky130_fd_sc_hd__buf_1 $T=83720 269280 0 0 $X=83530 $Y=269040
X1197 1 2 76 2 56 1 sky130_fd_sc_hd__buf_1 $T=103500 285600 0 0 $X=103310 $Y=285360
X1198 1 2 79 2 67 1 sky130_fd_sc_hd__buf_1 $T=105340 301920 1 0 $X=105150 $Y=298960
X1199 1 2 55 2 75 1 sky130_fd_sc_hd__buf_1 $T=106260 269280 0 0 $X=106070 $Y=269040
X1200 1 2 57 2 377 1 sky130_fd_sc_hd__buf_1 $T=111320 269280 0 0 $X=111130 $Y=269040
X1201 1 2 62 2 84 1 sky130_fd_sc_hd__buf_1 $T=115460 274720 1 0 $X=115270 $Y=271760
X1202 1 2 79 2 85 1 sky130_fd_sc_hd__buf_1 $T=116380 296480 1 0 $X=116190 $Y=293520
X1203 1 2 76 2 87 1 sky130_fd_sc_hd__buf_1 $T=119140 291040 0 0 $X=118950 $Y=290800
X1204 1 2 77 2 82 1 sky130_fd_sc_hd__buf_1 $T=119140 307360 0 0 $X=118950 $Y=307120
X1205 1 2 88 2 78 1 sky130_fd_sc_hd__buf_1 $T=120520 307360 1 0 $X=120330 $Y=304400
X1206 1 2 399 2 95 1 sky130_fd_sc_hd__buf_1 $T=151340 301920 1 0 $X=151150 $Y=298960
X1207 1 2 114 2 361 1 sky130_fd_sc_hd__buf_1 $T=151800 296480 1 0 $X=151610 $Y=293520
X1208 1 2 115 2 359 1 sky130_fd_sc_hd__buf_1 $T=151800 296480 0 0 $X=151610 $Y=296240
X1209 1 2 114 2 108 1 sky130_fd_sc_hd__buf_1 $T=153180 307360 0 0 $X=152990 $Y=307120
X1210 1 2 399 2 351 1 sky130_fd_sc_hd__buf_1 $T=155480 291040 0 0 $X=155290 $Y=290800
X1211 1 2 115 2 107 1 sky130_fd_sc_hd__buf_1 $T=158240 307360 0 0 $X=158050 $Y=307120
X1212 1 2 120 2 42 1 sky130_fd_sc_hd__buf_1 $T=159160 263840 0 0 $X=158970 $Y=263600
X1213 1 2 121 2 106 1 sky130_fd_sc_hd__buf_1 $T=161000 291040 0 0 $X=160810 $Y=290800
X1214 1 2 121 2 364 1 sky130_fd_sc_hd__buf_1 $T=162840 285600 1 0 $X=162650 $Y=282640
X1215 1 2 120 2 399 1 sky130_fd_sc_hd__buf_1 $T=168360 291040 1 0 $X=168170 $Y=288080
X1216 1 2 114 2 402 1 sky130_fd_sc_hd__buf_1 $T=168820 274720 0 0 $X=168630 $Y=274480
X1217 1 2 399 2 125 1 sky130_fd_sc_hd__buf_1 $T=168820 301920 0 0 $X=168630 $Y=301680
X1218 1 2 114 2 127 1 sky130_fd_sc_hd__buf_1 $T=169740 301920 1 0 $X=169550 $Y=298960
X1219 1 2 115 2 406 1 sky130_fd_sc_hd__buf_1 $T=175260 274720 0 0 $X=175070 $Y=274480
X1220 1 2 120 2 79 1 sky130_fd_sc_hd__buf_1 $T=175260 285600 0 0 $X=175070 $Y=285360
X1221 1 2 399 2 131 1 sky130_fd_sc_hd__buf_1 $T=176640 285600 1 0 $X=176450 $Y=282640
X1222 1 2 399 2 124 1 sky130_fd_sc_hd__buf_1 $T=179400 296480 1 0 $X=179210 $Y=293520
X1223 1 2 121 2 134 1 sky130_fd_sc_hd__buf_1 $T=189520 269280 1 0 $X=189330 $Y=266320
X1224 1 2 141 2 121 1 sky130_fd_sc_hd__buf_1 $T=192740 263840 0 0 $X=192550 $Y=263600
X1225 1 2 426 2 138 1 sky130_fd_sc_hd__buf_1 $T=203320 296480 0 0 $X=203130 $Y=296240
X1226 1 2 141 2 62 1 sky130_fd_sc_hd__buf_1 $T=207000 263840 0 0 $X=206810 $Y=263600
X1227 1 2 141 2 426 1 sky130_fd_sc_hd__buf_1 $T=209300 274720 1 0 $X=209110 $Y=271760
X1228 1 2 120 2 159 1 sky130_fd_sc_hd__buf_1 $T=212520 296480 0 0 $X=212330 $Y=296240
X1229 1 2 141 2 162 1 sky130_fd_sc_hd__buf_1 $T=217580 269280 1 0 $X=217390 $Y=266320
X1230 1 2 162 2 142 1 sky130_fd_sc_hd__buf_1 $T=220340 296480 0 0 $X=220150 $Y=296240
X1231 1 2 444 2 147 1 sky130_fd_sc_hd__buf_1 $T=226320 296480 1 0 $X=226130 $Y=293520
X1232 1 2 445 2 151 1 sky130_fd_sc_hd__buf_1 $T=231380 296480 1 0 $X=231190 $Y=293520
X1233 1 2 444 2 166 1 sky130_fd_sc_hd__buf_1 $T=234140 307360 1 0 $X=233950 $Y=304400
X1234 1 2 162 2 175 1 sky130_fd_sc_hd__buf_1 $T=237360 301920 0 0 $X=237170 $Y=301680
X1235 1 2 445 2 167 1 sky130_fd_sc_hd__buf_1 $T=239200 307360 1 0 $X=239010 $Y=304400
X1236 1 2 159 2 172 1 sky130_fd_sc_hd__buf_1 $T=241040 307360 0 0 $X=240850 $Y=307120
X1237 1 2 444 2 182 1 sky130_fd_sc_hd__buf_1 $T=253000 301920 0 0 $X=252810 $Y=301680
X1238 1 2 426 2 181 1 sky130_fd_sc_hd__buf_1 $T=259440 291040 0 0 $X=259250 $Y=290800
X1239 1 2 445 2 184 1 sky130_fd_sc_hd__buf_1 $T=267720 301920 0 0 $X=267530 $Y=301680
X1240 1 2 444 2 186 1 sky130_fd_sc_hd__buf_1 $T=272320 285600 0 0 $X=272130 $Y=285360
X1241 1 2 445 2 462 1 sky130_fd_sc_hd__buf_1 $T=273700 285600 1 0 $X=273510 $Y=282640
X1242 1 2 196 2 445 1 sky130_fd_sc_hd__buf_1 $T=278760 285600 1 0 $X=278570 $Y=282640
X1243 1 2 426 2 459 1 sky130_fd_sc_hd__buf_1 $T=280140 291040 0 0 $X=279950 $Y=290800
X1244 1 2 159 2 192 1 sky130_fd_sc_hd__buf_1 $T=280600 301920 0 0 $X=280410 $Y=301680
X1245 1 2 200 2 444 1 sky130_fd_sc_hd__buf_1 $T=283820 285600 1 0 $X=283630 $Y=282640
X1246 1 2 426 2 190 1 sky130_fd_sc_hd__buf_1 $T=284280 280160 1 0 $X=284090 $Y=277200
X1247 1 2 200 2 472 1 sky130_fd_sc_hd__buf_1 $T=292560 291040 1 0 $X=292370 $Y=288080
X1248 1 2 426 2 485 1 sky130_fd_sc_hd__buf_1 $T=295780 285600 0 0 $X=295590 $Y=285360
X1249 1 2 196 2 198 1 sky130_fd_sc_hd__buf_1 $T=296240 291040 0 0 $X=296050 $Y=290800
X1250 1 2 200 2 210 1 sky130_fd_sc_hd__buf_1 $T=298080 280160 0 0 $X=297890 $Y=279920
X1251 1 2 196 2 216 1 sky130_fd_sc_hd__buf_1 $T=302220 285600 0 0 $X=302030 $Y=285360
X1252 1 2 40 334 47 2 339 1 sky130_fd_sc_hd__o21a_4 $T=50140 269280 0 0 $X=49950 $Y=269040
X1253 1 2 48 328 45 2 338 1 sky130_fd_sc_hd__o21a_4 $T=50600 296480 1 0 $X=50410 $Y=293520
X1254 1 2 43 41 45 2 337 1 sky130_fd_sc_hd__o21a_4 $T=51980 301920 0 0 $X=51790 $Y=301680
X1255 1 2 44 331 45 2 344 1 sky130_fd_sc_hd__o21a_4 $T=52440 291040 0 0 $X=52250 $Y=290800
X1256 1 2 46 34 45 2 335 1 sky130_fd_sc_hd__o21a_4 $T=52440 307360 0 0 $X=52250 $Y=307120
X1257 1 2 50 343 47 2 341 1 sky130_fd_sc_hd__o21a_4 $T=54740 285600 1 0 $X=54550 $Y=282640
X1258 1 2 52 49 47 2 346 1 sky130_fd_sc_hd__o21a_4 $T=60720 280160 1 0 $X=60530 $Y=277200
X1259 1 2 59 61 47 2 348 1 sky130_fd_sc_hd__o21a_4 $T=63020 263840 0 0 $X=62830 $Y=263600
X1260 1 2 58 53 45 2 347 1 sky130_fd_sc_hd__o21a_4 $T=66700 307360 0 0 $X=66510 $Y=307120
X1261 1 2 63 350 47 2 354 1 sky130_fd_sc_hd__o21a_4 $T=72220 269280 0 0 $X=72030 $Y=269040
X1262 1 2 58 357 364 2 362 1 sky130_fd_sc_hd__o21a_4 $T=81420 296480 1 0 $X=81230 $Y=293520
X1263 1 2 43 368 364 2 370 1 sky130_fd_sc_hd__o21a_4 $T=88320 301920 1 0 $X=88130 $Y=298960
X1264 1 2 48 363 364 2 365 1 sky130_fd_sc_hd__o21a_4 $T=92460 291040 1 0 $X=92270 $Y=288080
X1265 1 2 80 372 84 2 376 1 sky130_fd_sc_hd__o21a_4 $T=106720 274720 0 0 $X=106530 $Y=274480
X1266 1 2 81 73 84 2 83 1 sky130_fd_sc_hd__o21a_4 $T=107180 263840 0 0 $X=106990 $Y=263600
X1267 1 2 81 86 87 2 374 1 sky130_fd_sc_hd__o21a_4 $T=108560 307360 1 0 $X=108370 $Y=304400
X1268 1 2 93 382 84 2 380 1 sky130_fd_sc_hd__o21a_4 $T=120060 280160 1 0 $X=119870 $Y=277200
X1269 1 2 80 381 87 2 383 1 sky130_fd_sc_hd__o21a_4 $T=121440 301920 1 0 $X=121250 $Y=298960
X1270 1 2 97 384 84 2 385 1 sky130_fd_sc_hd__o21a_4 $T=126500 263840 0 0 $X=126310 $Y=263600
X1271 1 2 44 390 106 2 393 1 sky130_fd_sc_hd__o21a_4 $T=136160 301920 1 0 $X=135970 $Y=298960
X1272 1 2 46 396 364 2 395 1 sky130_fd_sc_hd__o21a_4 $T=147200 291040 0 0 $X=147010 $Y=290800
X1273 1 2 111 112 118 2 116 1 sky130_fd_sc_hd__o21a_4 $T=151800 301920 0 0 $X=151610 $Y=301680
X1274 1 2 122 401 364 2 403 1 sky130_fd_sc_hd__o21a_4 $T=163300 280160 0 0 $X=163110 $Y=279920
X1275 1 2 111 410 118 2 412 1 sky130_fd_sc_hd__o21a_4 $T=176640 296480 0 0 $X=176450 $Y=296240
X1276 1 2 130 409 134 2 411 1 sky130_fd_sc_hd__o21a_4 $T=178940 269280 0 0 $X=178750 $Y=269040
X1277 1 2 93 132 138 2 135 1 sky130_fd_sc_hd__o21a_4 $T=185840 307360 0 0 $X=185650 $Y=307120
X1278 1 2 139 418 134 2 414 1 sky130_fd_sc_hd__o21a_4 $T=188600 269280 0 0 $X=188410 $Y=269040
X1279 1 2 80 422 138 2 416 1 sky130_fd_sc_hd__o21a_4 $T=189520 301920 0 0 $X=189330 $Y=301680
X1280 1 2 144 420 134 2 421 1 sky130_fd_sc_hd__o21a_4 $T=198720 274720 1 0 $X=198530 $Y=271760
X1281 1 2 80 425 142 2 428 1 sky130_fd_sc_hd__o21a_4 $T=202400 296480 1 0 $X=202210 $Y=293520
X1282 1 2 93 155 142 2 429 1 sky130_fd_sc_hd__o21a_4 $T=205160 307360 1 0 $X=204970 $Y=304400
X1283 1 2 111 431 118 2 430 1 sky130_fd_sc_hd__o21a_4 $T=205620 285600 0 0 $X=205430 $Y=285360
X1284 1 2 160 158 156 2 157 1 sky130_fd_sc_hd__o21a_4 $T=212060 263840 0 0 $X=211870 $Y=263600
X1285 1 2 161 433 142 2 435 1 sky130_fd_sc_hd__o21a_4 $T=217580 296480 1 0 $X=217390 $Y=293520
X1286 1 2 63 439 142 2 436 1 sky130_fd_sc_hd__o21a_4 $T=218500 301920 0 0 $X=218310 $Y=301680
X1287 1 2 180 451 459 2 450 1 sky130_fd_sc_hd__o21a_4 $T=253460 280160 1 0 $X=253270 $Y=277200
X1288 1 2 122 463 181 2 461 1 sky130_fd_sc_hd__o21a_4 $T=259440 285600 0 0 $X=259250 $Y=285360
X1289 1 2 43 452 181 2 455 1 sky130_fd_sc_hd__o21a_4 $T=259440 301920 0 0 $X=259250 $Y=301680
X1290 1 2 46 458 181 2 187 1 sky130_fd_sc_hd__o21a_4 $T=260360 301920 1 0 $X=260170 $Y=298960
X1291 1 2 130 188 190 2 464 1 sky130_fd_sc_hd__o21a_4 $T=268180 263840 0 0 $X=267990 $Y=263600
X1292 1 2 160 197 459 2 474 1 sky130_fd_sc_hd__o21a_4 $T=285200 301920 1 0 $X=285010 $Y=298960
X1293 1 2 139 473 190 2 469 1 sky130_fd_sc_hd__o21a_4 $T=287500 269280 0 0 $X=287310 $Y=269040
X1294 1 2 201 475 459 2 478 1 sky130_fd_sc_hd__o21a_4 $T=287500 285600 0 0 $X=287310 $Y=285360
X1295 1 2 144 479 190 2 476 1 sky130_fd_sc_hd__o21a_4 $T=290720 274720 0 0 $X=290530 $Y=274480
X1296 1 2 206 483 459 2 482 1 sky130_fd_sc_hd__o21a_4 $T=291640 296480 0 0 $X=291450 $Y=296240
X1297 1 2 213 211 485 2 486 1 sky130_fd_sc_hd__o21a_4 $T=301760 274720 1 0 $X=301570 $Y=271760
X1298 1 2 214 209 485 2 487 1 sky130_fd_sc_hd__o21a_4 $T=301760 301920 1 0 $X=301570 $Y=298960
X1299 1 2 218 494 190 2 491 1 sky130_fd_sc_hd__o21a_4 $T=304520 269280 0 0 $X=304330 $Y=269040
X1300 1 2 219 212 485 2 220 1 sky130_fd_sc_hd__o21a_4 $T=304980 301920 0 0 $X=304790 $Y=301680
X1301 1 2 222 489 459 2 488 1 sky130_fd_sc_hd__o21a_4 $T=305440 291040 1 0 $X=305250 $Y=288080
X1302 1 2 225 223 485 2 224 1 sky130_fd_sc_hd__o21a_4 $T=310040 301920 1 0 $X=309850 $Y=298960
X1303 1 2 226 227 485 2 499 1 sky130_fd_sc_hd__o21a_4 $T=315560 301920 0 0 $X=315370 $Y=301680
X1304 1 2 3 5 ICV_21 $T=18860 307360 0 0 $X=18670 $Y=307120
X1305 1 2 32 333 ICV_21 $T=38640 280160 1 0 $X=38450 $Y=277200
X1306 1 2 336 340 ICV_21 $T=43240 269280 0 0 $X=43050 $Y=269040
X1307 1 2 341 340 ICV_21 $T=45540 280160 0 0 $X=45350 $Y=279920
X1308 1 2 49 47 ICV_21 $T=54740 274720 0 0 $X=54550 $Y=274480
X1309 1 2 47 348 ICV_21 $T=70840 274720 1 0 $X=70650 $Y=271760
X1310 1 2 351 359 ICV_21 $T=74520 296480 0 0 $X=74330 $Y=296240
X1311 1 2 357 361 ICV_21 $T=76360 296480 1 0 $X=76170 $Y=293520
X1312 1 2 5 66 ICV_21 $T=81420 307360 0 0 $X=81230 $Y=307120
X1313 1 2 364 359 ICV_21 $T=86940 296480 1 0 $X=86750 $Y=293520
X1314 1 2 372 75 ICV_21 $T=99360 269280 0 0 $X=99170 $Y=269040
X1315 1 2 94 96 ICV_21 $T=121900 307360 1 0 $X=121710 $Y=304400
X1316 1 2 388 389 ICV_21 $T=125120 291040 1 0 $X=124930 $Y=288080
X1317 1 2 395 396 ICV_21 $T=138460 291040 1 0 $X=138270 $Y=288080
X1318 1 2 398 117 ICV_21 $T=148580 285600 1 0 $X=148390 $Y=282640
X1319 1 2 351 403 ICV_21 $T=159160 269280 0 0 $X=158970 $Y=269040
X1320 1 2 143 147 ICV_21 $T=196880 307360 0 0 $X=196690 $Y=307120
X1321 1 2 170 172 ICV_21 $T=230460 307360 0 0 $X=230270 $Y=307120
X1322 1 2 445 5 ICV_21 $T=241040 285600 0 0 $X=240850 $Y=285360
X1323 1 2 452 444 ICV_21 $T=247940 301920 0 0 $X=247750 $Y=301680
X1324 1 2 5 454 ICV_21 $T=249320 263840 0 0 $X=249130 $Y=263600
X1325 1 2 455 452 ICV_21 $T=250240 301920 1 0 $X=250050 $Y=298960
X1326 1 2 197 459 ICV_21 $T=281060 296480 0 0 $X=280870 $Y=296240
X1327 1 2 3 5 ICV_21 $T=333500 269280 0 0 $X=333310 $Y=269040
X1328 1 2 3 ICV_22 $T=6900 291040 0 0 $X=6710 $Y=290800
X1329 1 2 3 ICV_22 $T=6900 296480 0 0 $X=6710 $Y=296240
X1330 1 2 322 ICV_22 $T=34040 301920 0 0 $X=33850 $Y=301680
X1331 1 2 334 ICV_22 $T=48760 274720 0 0 $X=48570 $Y=274480
X1332 1 2 51 ICV_22 $T=57500 307360 1 0 $X=57310 $Y=304400
X1333 1 2 350 ICV_22 $T=66240 280160 1 0 $X=66050 $Y=277200
X1334 1 2 62 ICV_22 $T=67620 280160 0 0 $X=67430 $Y=279920
X1335 1 2 57 ICV_22 $T=68540 274720 1 0 $X=68350 $Y=271760
X1336 1 2 369 ICV_22 $T=86480 274720 0 0 $X=86290 $Y=274480
X1337 1 2 376 ICV_22 $T=100740 269280 1 0 $X=100550 $Y=266320
X1338 1 2 79 ICV_22 $T=103040 296480 0 0 $X=102850 $Y=296240
X1339 1 2 85 ICV_22 $T=105340 296480 0 0 $X=105150 $Y=296240
X1340 1 2 377 ICV_22 $T=118220 269280 0 0 $X=118030 $Y=269040
X1341 1 2 95 ICV_22 $T=122820 291040 1 0 $X=122630 $Y=288080
X1342 1 2 387 ICV_22 $T=124660 285600 1 0 $X=124470 $Y=282640
X1343 1 2 5 ICV_22 $T=142140 285600 0 0 $X=141950 $Y=285360
X1344 1 2 46 ICV_22 $T=142600 291040 0 0 $X=142410 $Y=290800
X1345 1 2 119 ICV_22 $T=151800 269280 0 0 $X=151610 $Y=269040
X1346 1 2 417 ICV_22 $T=181700 285600 1 0 $X=181510 $Y=282640
X1347 1 2 138 ICV_22 $T=184460 307360 1 0 $X=184270 $Y=304400
X1348 1 2 420 ICV_22 $T=184920 269280 1 0 $X=184730 $Y=266320
X1349 1 2 131 ICV_22 $T=192280 280160 1 0 $X=192090 $Y=277200
X1350 1 2 152 ICV_22 $T=202400 285600 0 0 $X=202210 $Y=285360
X1351 1 2 63 ICV_22 $T=215280 301920 0 0 $X=215090 $Y=301680
X1352 1 2 168 ICV_22 $T=224480 269280 0 0 $X=224290 $Y=269040
X1353 1 2 169 ICV_22 $T=226780 285600 0 0 $X=226590 $Y=285360
X1354 1 2 176 ICV_22 $T=237360 269280 1 0 $X=237170 $Y=266320
X1355 1 2 448 ICV_22 $T=238740 291040 1 0 $X=238550 $Y=288080
X1356 1 2 5 ICV_22 $T=265880 307360 0 0 $X=265690 $Y=307120
X1357 1 2 179 ICV_22 $T=273700 263840 0 0 $X=273510 $Y=263600
X1358 1 2 196 ICV_22 $T=277380 280160 0 0 $X=277190 $Y=279920
X1359 1 2 472 ICV_22 $T=277380 301920 0 0 $X=277190 $Y=301680
X1360 1 2 459 ICV_22 $T=285200 285600 1 0 $X=285010 $Y=282640
X1361 1 2 198 ICV_22 $T=286580 301920 0 0 $X=286390 $Y=301680
X1362 1 2 206 ICV_22 $T=288420 296480 0 0 $X=288230 $Y=296240
X1363 1 2 196 ICV_22 $T=299000 285600 0 0 $X=298810 $Y=285360
X1364 1 2 219 ICV_22 $T=301760 301920 0 0 $X=301570 $Y=301680
X1365 1 2 192 ICV_22 $T=303140 280160 0 0 $X=302950 $Y=279920
X1366 1 2 500 ICV_22 $T=314640 280160 0 0 $X=314450 $Y=279920
X1367 1 2 465 ICV_22 $T=328900 280160 1 0 $X=328710 $Y=277200
X1368 1 2 ICV_23 $T=20240 301920 1 0 $X=20050 $Y=298960
X1369 1 2 ICV_23 $T=20700 296480 0 0 $X=20510 $Y=296240
X1370 1 2 ICV_23 $T=34040 274720 0 0 $X=33850 $Y=274480
X1371 1 2 ICV_23 $T=76360 280160 1 0 $X=76170 $Y=277200
X1372 1 2 ICV_23 $T=76360 307360 1 0 $X=76170 $Y=304400
X1373 1 2 ICV_23 $T=91540 285600 1 0 $X=91350 $Y=282640
X1374 1 2 ICV_23 $T=104420 285600 1 0 $X=104230 $Y=282640
X1375 1 2 ICV_23 $T=118220 280160 0 0 $X=118030 $Y=279920
X1376 1 2 ICV_23 $T=132020 263840 0 0 $X=131830 $Y=263600
X1377 1 2 ICV_23 $T=137540 285600 1 0 $X=137350 $Y=282640
X1378 1 2 ICV_23 $T=138460 307360 1 0 $X=138270 $Y=304400
X1379 1 2 ICV_23 $T=139840 269280 1 0 $X=139650 $Y=266320
X1380 1 2 ICV_23 $T=154100 285600 0 0 $X=153910 $Y=285360
X1381 1 2 ICV_23 $T=168360 280160 1 0 $X=168170 $Y=277200
X1382 1 2 ICV_23 $T=169740 291040 1 0 $X=169550 $Y=288080
X1383 1 2 ICV_23 $T=186760 291040 0 0 $X=186570 $Y=290800
X1384 1 2 ICV_23 $T=188600 296480 1 0 $X=188410 $Y=293520
X1385 1 2 ICV_23 $T=207460 274720 0 0 $X=207270 $Y=274480
X1386 1 2 ICV_23 $T=213440 269280 0 0 $X=213250 $Y=269040
X1387 1 2 ICV_23 $T=227700 291040 1 0 $X=227510 $Y=288080
X1388 1 2 ICV_23 $T=230460 274720 0 0 $X=230270 $Y=274480
X1389 1 2 ICV_23 $T=236900 269280 0 0 $X=236710 $Y=269040
X1390 1 2 ICV_23 $T=236900 296480 0 0 $X=236710 $Y=296240
X1391 1 2 ICV_23 $T=244720 296480 1 0 $X=244530 $Y=293520
X1392 1 2 ICV_23 $T=258520 274720 0 0 $X=258330 $Y=274480
X1393 1 2 ICV_23 $T=270020 296480 0 0 $X=269830 $Y=296240
X1394 1 2 ICV_23 $T=287500 285600 1 0 $X=287310 $Y=282640
X1395 1 2 ICV_23 $T=312800 280160 1 0 $X=312610 $Y=277200
X1396 1 2 ICV_23 $T=316940 280160 0 0 $X=316750 $Y=279920
X1397 1 2 ICV_23 $T=319700 263840 0 0 $X=319510 $Y=263600
X1398 1 2 ICV_24 $T=18400 291040 1 0 $X=18210 $Y=288080
X1399 1 2 ICV_24 $T=18400 307360 1 0 $X=18210 $Y=304400
X1400 1 2 ICV_24 $T=74520 307360 1 0 $X=74330 $Y=304400
X1401 1 2 ICV_24 $T=102580 285600 1 0 $X=102390 $Y=282640
X1402 1 2 ICV_24 $T=116380 269280 0 0 $X=116190 $Y=269040
X1403 1 2 ICV_24 $T=116380 280160 0 0 $X=116190 $Y=279920
X1404 1 2 ICV_24 $T=116380 296480 0 0 $X=116190 $Y=296240
X1405 1 2 ICV_24 $T=130640 285600 1 0 $X=130450 $Y=282640
X1406 1 2 ICV_24 $T=130640 301920 1 0 $X=130450 $Y=298960
X1407 1 2 ICV_24 $T=144440 280160 0 0 $X=144250 $Y=279920
X1408 1 2 ICV_24 $T=144440 285600 0 0 $X=144250 $Y=285360
X1409 1 2 ICV_24 $T=158700 296480 1 0 $X=158510 $Y=293520
X1410 1 2 ICV_24 $T=186760 307360 1 0 $X=186570 $Y=304400
X1411 1 2 ICV_24 $T=242880 280160 1 0 $X=242690 $Y=277200
X1412 1 2 ICV_24 $T=312800 291040 0 0 $X=312610 $Y=290800
X1413 1 2 ICV_24 $T=312800 307360 0 0 $X=312610 $Y=307120
.ENDS
***************************************
.SUBCKT ICV_26 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 5440 1 0 $X=-190 $Y=2480
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3
** N=3 EP=3 IP=5 FDC=3
*.SEEDPROM
X1 1 2 3 ICV_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_29 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=17
*.SEEDPROM
X0 1 3 sky130_fd_sc_hd__diode_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 4 5 2 6 1 sky130_fd_sc_hd__nor2_4 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254
** N=591 EP=254 IP=5655 FDC=8601
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=221625 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=227065 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=232505 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=237945 $D=191
X4 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=243385 $D=191
X5 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=248825 $D=191
X6 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=254265 $D=191
X7 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=259705 $D=191
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 220320 1 0 $X=5330 $Y=217360
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28060 231200 1 0 $X=27870 $Y=228240
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=37260 236640 1 0 $X=37070 $Y=233680
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=38640 263840 1 0 $X=38450 $Y=260880
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=56120 263840 1 0 $X=55930 $Y=260880
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=65320 225760 1 0 $X=65130 $Y=222800
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74980 225760 0 0 $X=74790 $Y=225520
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 220320 1 0 $X=76170 $Y=217360
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 247520 1 0 $X=76170 $Y=244560
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 220320 1 0 $X=102390 $Y=217360
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=117300 263840 1 0 $X=117110 $Y=260880
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=117760 231200 1 0 $X=117570 $Y=228240
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=122360 258400 1 0 $X=122170 $Y=255440
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=149960 236640 1 0 $X=149770 $Y=233680
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=150880 225760 1 0 $X=150690 $Y=222800
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 220320 1 0 $X=158510 $Y=217360
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174800 263840 1 0 $X=174610 $Y=260880
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=200560 220320 1 0 $X=200370 $Y=217360
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=222180 220320 1 0 $X=221990 $Y=217360
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 225760 0 0 $X=230270 $Y=225520
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=237360 242080 1 0 $X=237170 $Y=239120
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=257140 220320 1 0 $X=256950 $Y=217360
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=257140 231200 1 0 $X=256950 $Y=228240
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=274620 231200 0 0 $X=274430 $Y=230960
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=283820 263840 1 0 $X=283630 $Y=260880
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=293940 225760 0 0 $X=293750 $Y=225520
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=306820 220320 1 0 $X=306630 $Y=217360
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=310040 252960 1 0 $X=309850 $Y=250000
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=327060 225760 1 0 $X=326870 $Y=222800
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 247520 0 0 $X=340670 $Y=247280
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 252960 0 0 $X=340670 $Y=252720
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 220320 0 180 $X=348950 $Y=217360
X143 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=10580 225760 1 0 $X=10390 $Y=222800
X144 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 225760 1 0 $X=20050 $Y=222800
X145 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 247520 1 0 $X=20050 $Y=244560
X146 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=42780 242080 1 0 $X=42590 $Y=239120
X147 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 236640 1 0 $X=43970 $Y=233680
X148 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 247520 1 0 $X=43970 $Y=244560
X149 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 258400 1 0 $X=43970 $Y=255440
X150 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=48300 258400 1 0 $X=48110 $Y=255440
X151 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=59340 231200 1 0 $X=59150 $Y=228240
X152 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=61640 225760 1 0 $X=61450 $Y=222800
X153 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=62100 252960 0 0 $X=61910 $Y=252720
X154 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=64400 252960 1 0 $X=64210 $Y=250000
X155 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=66700 236640 1 0 $X=66510 $Y=233680
X156 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=70840 258400 1 0 $X=70650 $Y=255440
X157 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 252960 1 0 $X=72030 $Y=250000
X158 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=86020 247520 0 0 $X=85830 $Y=247280
X159 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=91540 242080 1 0 $X=91350 $Y=239120
X160 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=95680 252960 0 0 $X=95490 $Y=252720
X161 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=98900 220320 1 0 $X=98710 $Y=217360
X162 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=98900 225760 1 0 $X=98710 $Y=222800
X163 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 236640 1 0 $X=100090 $Y=233680
X164 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 236640 1 0 $X=104230 $Y=233680
X165 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 242080 1 0 $X=104230 $Y=239120
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=114080 231200 1 0 $X=113890 $Y=228240
X167 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=116380 220320 1 0 $X=116190 $Y=217360
X168 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=118220 231200 0 0 $X=118030 $Y=230960
X169 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126500 220320 1 0 $X=126310 $Y=217360
X170 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 247520 1 0 $X=132290 $Y=244560
X171 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=138920 236640 1 0 $X=138730 $Y=233680
X172 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=141680 220320 0 0 $X=141490 $Y=220080
X173 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 220320 0 0 $X=146090 $Y=220080
X174 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=148580 220320 1 0 $X=148390 $Y=217360
X175 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 231200 1 0 $X=156210 $Y=228240
X176 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=163300 247520 0 0 $X=163110 $Y=247280
X177 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=164220 252960 1 0 $X=164030 $Y=250000
X178 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=167900 242080 1 0 $X=167710 $Y=239120
X179 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=171120 263840 1 0 $X=170930 $Y=260880
X180 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=177100 252960 1 0 $X=176910 $Y=250000
X181 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183540 242080 1 0 $X=183350 $Y=239120
X182 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183540 263840 1 0 $X=183350 $Y=260880
X183 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 247520 1 0 $X=184270 $Y=244560
X184 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198260 258400 0 0 $X=198070 $Y=258160
X185 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=203320 220320 1 0 $X=203130 $Y=217360
X186 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=204240 225760 1 0 $X=204050 $Y=222800
X187 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212060 225760 1 0 $X=211870 $Y=222800
X188 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 252960 1 0 $X=212330 $Y=250000
X189 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 236640 0 0 $X=216470 $Y=236400
X190 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=221260 225760 0 0 $X=221070 $Y=225520
X191 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=227700 236640 1 0 $X=227510 $Y=233680
X192 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 252960 0 0 $X=230270 $Y=252720
X193 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239200 220320 0 0 $X=239010 $Y=220080
X194 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240120 242080 1 0 $X=239930 $Y=239120
X195 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 225760 1 0 $X=240390 $Y=222800
X196 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=241960 247520 0 0 $X=241770 $Y=247280
X197 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249780 263840 1 0 $X=249590 $Y=260880
X198 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254380 258400 1 0 $X=254190 $Y=255440
X199 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258520 258400 0 0 $X=258330 $Y=258160
X200 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=263580 231200 0 0 $X=263390 $Y=230960
X201 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=265880 220320 0 0 $X=265690 $Y=220080
X202 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267260 225760 1 0 $X=267070 $Y=222800
X203 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 252960 1 0 $X=268450 $Y=250000
X204 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 258400 1 0 $X=268450 $Y=255440
X205 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 242080 1 0 $X=272590 $Y=239120
X206 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281520 225760 1 0 $X=281330 $Y=222800
X207 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 231200 1 0 $X=296510 $Y=228240
X208 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 258400 1 0 $X=296510 $Y=255440
X209 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=297620 247520 0 0 $X=297430 $Y=247280
X210 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=299000 252960 0 0 $X=298810 $Y=252720
X211 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 247520 1 0 $X=300650 $Y=244560
X212 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 252960 1 0 $X=300650 $Y=250000
X213 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 258400 1 0 $X=300650 $Y=255440
X214 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=301760 258400 0 0 $X=301570 $Y=258160
X215 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=306820 242080 1 0 $X=306630 $Y=239120
X216 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=306820 247520 1 0 $X=306630 $Y=244560
X217 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 242080 1 0 $X=324570 $Y=239120
X218 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=330740 225760 0 0 $X=330550 $Y=225520
X219 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=331200 231200 1 0 $X=331010 $Y=228240
X220 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 252960 1 0 $X=344810 $Y=250000
X221 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 220320 1 0 $X=345270 $Y=217360
X222 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 225760 1 0 $X=345270 $Y=222800
X223 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 231200 1 0 $X=345270 $Y=228240
X224 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 242080 1 0 $X=345270 $Y=239120
X225 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 247520 1 0 $X=345270 $Y=244560
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 263840 1 0 $X=345270 $Y=260880
X227 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 225760 0 0 $X=6710 $Y=225520
X228 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 263840 1 0 $X=6710 $Y=260880
X229 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=28060 247520 0 0 $X=27870 $Y=247280
X230 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=28520 263840 1 0 $X=28330 $Y=260880
X231 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=39100 225760 1 0 $X=38910 $Y=222800
X232 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=41400 231200 1 0 $X=41210 $Y=228240
X233 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=45080 258400 0 0 $X=44890 $Y=258160
X234 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=53360 242080 1 0 $X=53170 $Y=239120
X235 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=54280 242080 0 0 $X=54090 $Y=241840
X236 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=64860 231200 1 0 $X=64670 $Y=228240
X237 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=68080 263840 1 0 $X=67890 $Y=260880
X238 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=73600 247520 0 0 $X=73410 $Y=247280
X239 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=76820 258400 0 0 $X=76630 $Y=258160
X240 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=84180 252960 0 0 $X=83990 $Y=252720
X241 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=87400 252960 1 0 $X=87210 $Y=250000
X242 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97060 258400 1 0 $X=96870 $Y=255440
X243 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=98440 231200 1 0 $X=98250 $Y=228240
X244 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=107180 242080 0 0 $X=106990 $Y=241840
X245 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=108100 247520 1 0 $X=107910 $Y=244560
X246 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=109940 247520 0 0 $X=109750 $Y=247280
X247 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=111780 252960 1 0 $X=111590 $Y=250000
X248 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=117760 225760 1 0 $X=117570 $Y=222800
X249 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=122820 242080 1 0 $X=122630 $Y=239120
X250 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=124200 247520 1 0 $X=124010 $Y=244560
X251 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=124200 252960 1 0 $X=124010 $Y=250000
X252 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 242080 0 0 $X=125390 $Y=241840
X253 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=126040 225760 1 0 $X=125850 $Y=222800
X254 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=137540 225760 1 0 $X=137350 $Y=222800
X255 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=142600 247520 1 0 $X=142410 $Y=244560
X256 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=143520 231200 1 0 $X=143330 $Y=228240
X257 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=143520 252960 1 0 $X=143330 $Y=250000
X258 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=149960 263840 1 0 $X=149770 $Y=260880
X259 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=154100 247520 0 0 $X=153910 $Y=247280
X260 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=182160 258400 1 0 $X=181970 $Y=255440
X261 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=193200 236640 0 0 $X=193010 $Y=236400
X262 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=194580 242080 0 0 $X=194390 $Y=241840
X263 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195960 225760 1 0 $X=195770 $Y=222800
X264 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195960 247520 1 0 $X=195770 $Y=244560
X265 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=224020 236640 0 0 $X=223830 $Y=236400
X266 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=230460 252960 1 0 $X=230270 $Y=250000
X267 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=231840 242080 1 0 $X=231650 $Y=239120
X268 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235520 242080 0 0 $X=235330 $Y=241840
X269 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235980 225760 0 0 $X=235790 $Y=225520
X270 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=236440 231200 1 0 $X=236250 $Y=228240
X271 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237360 220320 1 0 $X=237170 $Y=217360
X272 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=238280 263840 1 0 $X=238090 $Y=260880
X273 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=252080 252960 1 0 $X=251890 $Y=250000
X274 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=258980 263840 1 0 $X=258790 $Y=260880
X275 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=264040 220320 1 0 $X=263850 $Y=217360
X276 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=268640 258400 0 0 $X=268450 $Y=258160
X277 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=280600 242080 1 0 $X=280410 $Y=239120
X278 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293020 236640 1 0 $X=292830 $Y=233680
X279 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293480 225760 1 0 $X=293290 $Y=222800
X280 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=294860 247520 1 0 $X=294670 $Y=244560
X281 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=299920 242080 0 0 $X=299730 $Y=241840
X282 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=334420 231200 0 0 $X=334230 $Y=230960
X283 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=335340 247520 0 0 $X=335150 $Y=247280
X284 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=340400 236640 1 0 $X=340210 $Y=233680
X285 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=341320 258400 1 0 $X=341130 $Y=255440
X286 1 2 ICV_2 $T=33580 247520 0 0 $X=33390 $Y=247280
X287 1 2 ICV_2 $T=103960 220320 1 0 $X=103770 $Y=217360
X288 1 2 ICV_2 $T=103960 231200 1 0 $X=103770 $Y=228240
X289 1 2 ICV_2 $T=160080 220320 1 0 $X=159890 $Y=217360
X290 1 2 ICV_2 $T=216200 220320 1 0 $X=216010 $Y=217360
X291 1 2 ICV_2 $T=216200 225760 1 0 $X=216010 $Y=222800
X292 1 2 ICV_2 $T=230000 236640 0 0 $X=229810 $Y=236400
X293 1 2 ICV_2 $T=286120 242080 0 0 $X=285930 $Y=241840
X294 1 2 ICV_2 $T=300380 231200 1 0 $X=300190 $Y=228240
X295 1 2 ICV_2 $T=300380 236640 1 0 $X=300190 $Y=233680
X296 1 2 ICV_2 $T=328440 220320 1 0 $X=328250 $Y=217360
X297 1 2 ICV_2 $T=328440 225760 1 0 $X=328250 $Y=222800
X298 1 2 ICV_2 $T=328440 242080 1 0 $X=328250 $Y=239120
X299 1 2 ICV_2 $T=328440 247520 1 0 $X=328250 $Y=244560
X300 1 2 ICV_2 $T=328440 263840 1 0 $X=328250 $Y=260880
X301 1 2 ICV_2 $T=342240 220320 0 0 $X=342050 $Y=220080
X302 1 2 ICV_2 $T=342240 225760 0 0 $X=342050 $Y=225520
X303 1 2 ICV_2 $T=342240 231200 0 0 $X=342050 $Y=230960
X304 1 2 ICV_2 $T=342240 236640 0 0 $X=342050 $Y=236400
X305 1 2 ICV_2 $T=342240 242080 0 0 $X=342050 $Y=241840
X306 1 2 ICV_2 $T=342240 247520 0 0 $X=342050 $Y=247280
X307 1 2 ICV_2 $T=342240 252960 0 0 $X=342050 $Y=252720
X308 1 2 ICV_2 $T=342240 258400 0 0 $X=342050 $Y=258160
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 236640 1 0 $X=17750 $Y=233680
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 247520 0 0 $X=18210 $Y=247280
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=25300 225760 0 0 $X=25110 $Y=225520
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=29440 252960 0 0 $X=29250 $Y=252720
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=30360 247520 1 0 $X=30170 $Y=244560
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31280 258400 1 0 $X=31090 $Y=255440
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=32200 242080 1 0 $X=32010 $Y=239120
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 252960 0 0 $X=33850 $Y=252720
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46460 242080 0 0 $X=46270 $Y=241840
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=58880 242080 1 0 $X=58690 $Y=239120
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59800 242080 0 0 $X=59610 $Y=241840
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69000 220320 1 0 $X=68810 $Y=217360
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73600 263840 1 0 $X=73410 $Y=260880
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=92920 252960 1 0 $X=92730 $Y=250000
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=101660 242080 1 0 $X=101470 $Y=239120
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 236640 0 0 $X=104230 $Y=236400
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 247520 0 0 $X=118030 $Y=247280
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=123280 231200 1 0 $X=123090 $Y=228240
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=124200 263840 1 0 $X=124010 $Y=260880
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=130180 258400 1 0 $X=129990 $Y=255440
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=132940 258400 0 0 $X=132750 $Y=258160
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=153640 258400 0 0 $X=153450 $Y=258160
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=154100 252960 0 0 $X=153910 $Y=252720
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=155940 252960 1 0 $X=155750 $Y=250000
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172500 231200 1 0 $X=172310 $Y=228240
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=175720 242080 1 0 $X=175530 $Y=239120
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=178020 247520 1 0 $X=177830 $Y=244560
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188600 220320 1 0 $X=188410 $Y=217360
X337 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=191820 252960 0 0 $X=191630 $Y=252720
X338 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=199640 236640 1 0 $X=199450 $Y=233680
X339 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=200100 242080 0 0 $X=199910 $Y=241840
X340 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=200100 252960 0 0 $X=199910 $Y=252720
X341 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 247520 1 0 $X=216470 $Y=244560
X342 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=218960 252960 1 0 $X=218770 $Y=250000
X343 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=232760 231200 0 0 $X=232570 $Y=230960
X344 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=241500 225760 0 0 $X=241310 $Y=225520
X345 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=241960 231200 1 0 $X=241770 $Y=228240
X346 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 247520 1 0 $X=242230 $Y=244560
X347 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=245640 242080 0 0 $X=245450 $Y=241840
X348 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=281980 258400 0 0 $X=281790 $Y=258160
X349 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284740 231200 1 0 $X=284550 $Y=228240
X350 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286120 252960 1 0 $X=285930 $Y=250000
X351 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298080 242080 1 0 $X=297890 $Y=239120
X352 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 236640 1 0 $X=298350 $Y=233680
X353 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 220320 0 0 $X=325950 $Y=220080
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=339940 231200 0 0 $X=339750 $Y=230960
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=346840 258400 1 0 $X=346650 $Y=255440
X356 1 4 sky130_fd_sc_hd__diode_2 $T=12880 225760 0 0 $X=12690 $Y=225520
X357 1 351 sky130_fd_sc_hd__diode_2 $T=19320 242080 0 0 $X=19130 $Y=241840
X358 1 366 sky130_fd_sc_hd__diode_2 $T=34500 242080 1 0 $X=34310 $Y=239120
X359 1 30 sky130_fd_sc_hd__diode_2 $T=34960 236640 0 0 $X=34770 $Y=236400
X360 1 4 sky130_fd_sc_hd__diode_2 $T=38640 220320 0 0 $X=38450 $Y=220080
X361 1 35 sky130_fd_sc_hd__diode_2 $T=48760 231200 0 0 $X=48570 $Y=230960
X362 1 70 sky130_fd_sc_hd__diode_2 $T=80040 247520 0 0 $X=79850 $Y=247280
X363 1 389 sky130_fd_sc_hd__diode_2 $T=83720 231200 1 0 $X=83530 $Y=228240
X364 1 80 sky130_fd_sc_hd__diode_2 $T=102580 258400 0 0 $X=102390 $Y=258160
X365 1 97 sky130_fd_sc_hd__diode_2 $T=119140 225760 0 0 $X=118950 $Y=225520
X366 1 99 sky130_fd_sc_hd__diode_2 $T=120520 220320 0 0 $X=120330 $Y=220080
X367 1 425 sky130_fd_sc_hd__diode_2 $T=147200 242080 0 0 $X=147010 $Y=241840
X368 1 4 sky130_fd_sc_hd__diode_2 $T=150420 220320 0 0 $X=150230 $Y=220080
X369 1 4 sky130_fd_sc_hd__diode_2 $T=156400 252960 0 0 $X=156210 $Y=252720
X370 1 124 sky130_fd_sc_hd__diode_2 $T=158700 225760 0 0 $X=158510 $Y=225520
X371 1 134 sky130_fd_sc_hd__diode_2 $T=171120 236640 1 0 $X=170930 $Y=233680
X372 1 4 sky130_fd_sc_hd__diode_2 $T=179400 247520 0 0 $X=179210 $Y=247280
X373 1 156 sky130_fd_sc_hd__diode_2 $T=191820 258400 1 0 $X=191630 $Y=255440
X374 1 122 sky130_fd_sc_hd__diode_2 $T=205160 252960 1 0 $X=204970 $Y=250000
X375 1 472 sky130_fd_sc_hd__diode_2 $T=219420 242080 1 0 $X=219230 $Y=239120
X376 1 475 sky130_fd_sc_hd__diode_2 $T=222180 225760 1 0 $X=221990 $Y=222800
X377 1 184 sky130_fd_sc_hd__diode_2 $T=234140 252960 0 0 $X=233950 $Y=252720
X378 1 4 sky130_fd_sc_hd__diode_2 $T=235060 231200 0 0 $X=234870 $Y=230960
X379 1 187 sky130_fd_sc_hd__diode_2 $T=242880 258400 0 0 $X=242690 $Y=258160
X380 1 199 sky130_fd_sc_hd__diode_2 $T=260820 252960 0 0 $X=260630 $Y=252720
X381 1 4 sky130_fd_sc_hd__diode_2 $T=268180 236640 0 0 $X=267990 $Y=236400
X382 1 203 sky130_fd_sc_hd__diode_2 $T=273240 220320 0 0 $X=273050 $Y=220080
X383 1 209 sky130_fd_sc_hd__diode_2 $T=275080 263840 1 0 $X=274890 $Y=260880
X384 1 4 sky130_fd_sc_hd__diode_2 $T=280140 252960 1 0 $X=279950 $Y=250000
X385 1 192 sky130_fd_sc_hd__diode_2 $T=303140 252960 0 0 $X=302950 $Y=252720
X386 1 525 sky130_fd_sc_hd__diode_2 $T=304980 258400 1 0 $X=304790 $Y=255440
X387 1 526 sky130_fd_sc_hd__diode_2 $T=318320 242080 0 0 $X=318130 $Y=241840
X388 1 159 sky130_fd_sc_hd__diode_2 $T=318780 220320 0 0 $X=318590 $Y=220080
X389 1 199 sky130_fd_sc_hd__diode_2 $T=320620 236640 0 0 $X=320430 $Y=236400
X390 1 4 sky130_fd_sc_hd__diode_2 $T=323840 258400 0 0 $X=323650 $Y=258160
X391 1 242 sky130_fd_sc_hd__diode_2 $T=328440 220320 0 0 $X=328250 $Y=220080
X392 1 2 15 ICV_4 $T=23000 236640 0 0 $X=22810 $Y=236400
X393 1 2 23 ICV_4 $T=35880 231200 1 0 $X=35690 $Y=228240
X394 1 2 371 ICV_4 $T=48760 242080 0 0 $X=48570 $Y=241840
X395 1 2 41 ICV_4 $T=52900 258400 1 0 $X=52710 $Y=255440
X396 1 2 378 ICV_4 $T=63020 247520 1 0 $X=62830 $Y=244560
X397 1 2 383 ICV_4 $T=70840 231200 1 0 $X=70650 $Y=228240
X398 1 2 64 ICV_4 $T=71300 236640 1 0 $X=71110 $Y=233680
X399 1 2 48 ICV_4 $T=76360 225760 0 0 $X=76170 $Y=225520
X400 1 2 379 ICV_4 $T=78660 220320 0 0 $X=78470 $Y=220080
X401 1 2 68 ICV_4 $T=85560 225760 1 0 $X=85370 $Y=222800
X402 1 2 392 ICV_4 $T=89240 220320 1 0 $X=89050 $Y=217360
X403 1 2 72 ICV_4 $T=90160 258400 1 0 $X=89970 $Y=255440
X404 1 2 78 ICV_4 $T=96600 247520 0 0 $X=96410 $Y=247280
X405 1 2 90 ICV_4 $T=115000 220320 0 0 $X=114810 $Y=220080
X406 1 2 103 ICV_4 $T=128800 220320 0 0 $X=128610 $Y=220080
X407 1 2 119 ICV_4 $T=147200 258400 1 0 $X=147010 $Y=255440
X408 1 2 127 ICV_4 $T=165600 242080 0 0 $X=165410 $Y=241840
X409 1 2 440 ICV_4 $T=172960 252960 1 0 $X=172770 $Y=250000
X410 1 2 4 ICV_4 $T=176180 258400 1 0 $X=175990 $Y=255440
X411 1 2 447 ICV_4 $T=176180 263840 1 0 $X=175990 $Y=260880
X412 1 2 137 ICV_4 $T=177560 242080 0 0 $X=177370 $Y=241840
X413 1 2 134 ICV_4 $T=183080 231200 1 0 $X=182890 $Y=228240
X414 1 2 455 ICV_4 $T=183540 225760 1 0 $X=183350 $Y=222800
X415 1 2 449 ICV_4 $T=188600 231200 0 0 $X=188410 $Y=230960
X416 1 2 153 ICV_4 $T=193660 231200 0 0 $X=193470 $Y=230960
X417 1 2 158 ICV_4 $T=198720 231200 0 0 $X=198530 $Y=230960
X418 1 2 460 ICV_4 $T=202400 247520 1 0 $X=202210 $Y=244560
X419 1 2 138 ICV_4 $T=212980 231200 1 0 $X=212790 $Y=228240
X420 1 2 470 ICV_4 $T=212980 236640 1 0 $X=212790 $Y=233680
X421 1 2 465 ICV_4 $T=212980 258400 1 0 $X=212790 $Y=255440
X422 1 2 163 ICV_4 $T=213440 220320 1 0 $X=213250 $Y=217360
X423 1 2 177 ICV_4 $T=233680 220320 0 0 $X=233490 $Y=220080
X424 1 2 182 ICV_4 $T=234140 236640 1 0 $X=233950 $Y=233680
X425 1 2 480 ICV_4 $T=236440 252960 1 0 $X=236250 $Y=250000
X426 1 2 146 ICV_4 $T=238280 252960 0 0 $X=238090 $Y=252720
X427 1 2 490 ICV_4 $T=245640 220320 1 0 $X=245450 $Y=217360
X428 1 2 184 ICV_4 $T=247480 242080 0 0 $X=247290 $Y=241840
X429 1 2 481 ICV_4 $T=250240 247520 0 0 $X=250050 $Y=247280
X430 1 2 496 ICV_4 $T=255760 225760 1 0 $X=255570 $Y=222800
X431 1 2 488 ICV_4 $T=258520 231200 1 0 $X=258330 $Y=228240
X432 1 2 506 ICV_4 $T=273700 258400 1 0 $X=273510 $Y=255440
X433 1 2 203 ICV_4 $T=276000 231200 1 0 $X=275810 $Y=228240
X434 1 2 140 ICV_4 $T=278760 220320 1 0 $X=278570 $Y=217360
X435 1 2 513 ICV_4 $T=278760 236640 1 0 $X=278570 $Y=233680
X436 1 2 211 ICV_4 $T=281520 236640 0 0 $X=281330 $Y=236400
X437 1 2 145 ICV_4 $T=282900 225760 0 0 $X=282710 $Y=225520
X438 1 2 505 ICV_4 $T=283360 252960 0 0 $X=283170 $Y=252720
X439 1 2 224 ICV_4 $T=294860 220320 0 0 $X=294670 $Y=220080
X440 1 2 131 ICV_4 $T=304520 247520 0 0 $X=304330 $Y=247280
X441 1 2 141 ICV_4 $T=306820 263840 1 0 $X=306630 $Y=260880
X442 1 2 529 ICV_4 $T=308200 225760 1 0 $X=308010 $Y=222800
X443 1 2 198 ICV_4 $T=309580 258400 0 0 $X=309390 $Y=258160
X444 1 2 231 ICV_4 $T=315560 220320 0 0 $X=315370 $Y=220080
X445 1 2 448 ICV_4 $T=315560 242080 0 0 $X=315370 $Y=241840
X446 1 2 431 ICV_4 $T=316480 258400 1 0 $X=316290 $Y=255440
X447 1 2 532 ICV_4 $T=320620 258400 0 0 $X=320430 $Y=258160
X448 1 2 246 ICV_4 $T=339020 220320 0 0 $X=338830 $Y=220080
X449 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 258400 0 0 $X=6710 $Y=258160
X450 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=10580 258400 1 0 $X=10390 $Y=255440
X451 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=18400 220320 0 0 $X=18210 $Y=220080
X452 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=20240 220320 1 0 $X=20050 $Y=217360
X453 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=25300 242080 0 0 $X=25110 $Y=241840
X454 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=44620 225760 1 0 $X=44430 $Y=222800
X455 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 247520 1 0 $X=48110 $Y=244560
X456 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 263840 1 0 $X=48110 $Y=260880
X457 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=52440 225760 0 0 $X=52250 $Y=225520
X458 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=87400 258400 1 0 $X=87210 $Y=255440
X459 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 242080 0 0 $X=89970 $Y=241840
X460 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 247520 0 0 $X=89970 $Y=247280
X461 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 252960 0 0 $X=89970 $Y=252720
X462 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=108560 252960 0 0 $X=108370 $Y=252720
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=109940 231200 1 0 $X=109750 $Y=228240
X464 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=114540 252960 0 0 $X=114350 $Y=252720
X465 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 231200 0 0 $X=114810 $Y=230960
X466 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 242080 0 0 $X=114810 $Y=241840
X467 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=122820 236640 1 0 $X=122630 $Y=233680
X468 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=124660 236640 0 0 $X=124470 $Y=236400
X469 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=131100 242080 0 0 $X=130910 $Y=241840
X470 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 263840 1 0 $X=132290 $Y=260880
X471 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=137540 258400 1 0 $X=137350 $Y=255440
X472 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 225760 1 0 $X=142870 $Y=222800
X473 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 252960 0 0 $X=142870 $Y=252720
X474 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=144440 258400 1 0 $X=144250 $Y=255440
X475 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 231200 0 0 $X=146090 $Y=230960
X476 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 252960 0 0 $X=146090 $Y=252720
X477 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=149040 231200 1 0 $X=148850 $Y=228240
X478 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=166060 220320 1 0 $X=165870 $Y=217360
X479 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=166980 258400 1 0 $X=166790 $Y=255440
X480 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=166980 263840 1 0 $X=166790 $Y=260880
X481 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=167900 236640 1 0 $X=167710 $Y=233680
X482 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=171580 225760 1 0 $X=171390 $Y=222800
X483 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=176640 247520 0 0 $X=176450 $Y=247280
X484 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=183540 220320 1 0 $X=183350 $Y=217360
X485 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=184000 252960 0 0 $X=183810 $Y=252720
X486 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=198720 236640 0 0 $X=198530 $Y=236400
X487 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 252960 0 0 $X=202210 $Y=252720
X488 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 258400 0 0 $X=202210 $Y=258160
X489 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=206080 258400 1 0 $X=205890 $Y=255440
X490 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213900 242080 0 0 $X=213710 $Y=241840
X491 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 242080 1 0 $X=216470 $Y=239120
X492 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=223560 252960 1 0 $X=223370 $Y=250000
X493 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 252960 0 0 $X=226590 $Y=252720
X494 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=227700 258400 1 0 $X=227510 $Y=255440
X495 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=235980 236640 0 0 $X=235790 $Y=236400
X496 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 258400 1 0 $X=244530 $Y=255440
X497 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=254840 252960 0 0 $X=254650 $Y=252720
X498 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=267260 236640 1 0 $X=267070 $Y=233680
X499 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=278300 263840 1 0 $X=278110 $Y=260880
X500 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=283360 242080 0 0 $X=283170 $Y=241840
X501 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=345920 236640 1 0 $X=345730 $Y=233680
X502 1 2 4 ICV_5 $T=7820 236640 1 0 $X=7630 $Y=233680
X503 1 2 28 ICV_5 $T=34960 220320 0 0 $X=34770 $Y=220080
X504 1 2 35 ICV_5 $T=41400 231200 0 0 $X=41210 $Y=230960
X505 1 2 35 ICV_5 $T=57960 225760 0 0 $X=57770 $Y=225520
X506 1 2 382 ICV_5 $T=72220 242080 1 0 $X=72030 $Y=239120
X507 1 2 388 ICV_5 $T=96140 225760 0 0 $X=95950 $Y=225520
X508 1 2 132 ICV_5 $T=170200 258400 0 0 $X=170010 $Y=258160
X509 1 2 136 ICV_5 $T=174800 225760 1 0 $X=174610 $Y=222800
X510 1 2 453 ICV_5 $T=198260 220320 0 0 $X=198070 $Y=220080
X511 1 2 183 ICV_5 $T=232760 225760 1 0 $X=232570 $Y=222800
X512 1 2 503 ICV_5 $T=264500 263840 1 0 $X=264310 $Y=260880
X513 1 2 201 ICV_5 $T=268180 263840 1 0 $X=267990 $Y=260880
X514 1 2 508 ICV_5 $T=268640 247520 1 0 $X=268450 $Y=244560
X515 1 2 214 ICV_5 $T=281980 247520 0 0 $X=281790 $Y=247280
X516 1 2 4 ICV_5 $T=288420 252960 1 0 $X=288230 $Y=250000
X517 1 2 221 ICV_5 $T=288420 258400 1 0 $X=288230 $Y=255440
X518 1 2 137 ICV_5 $T=305440 242080 0 0 $X=305250 $Y=241840
X519 1 2 539 ICV_5 $T=324300 236640 1 0 $X=324110 $Y=233680
X520 1 2 247 ICV_5 $T=338560 225760 0 0 $X=338370 $Y=225520
X521 1 2 541 ICV_5 $T=338560 236640 0 0 $X=338370 $Y=236400
X522 1 2 248 ICV_5 $T=338560 242080 0 0 $X=338370 $Y=241840
X523 1 2 354 ICV_6 $T=14720 225760 1 0 $X=14530 $Y=222800
X524 1 2 21 ICV_6 $T=28060 220320 0 0 $X=27870 $Y=220080
X525 1 2 29 ICV_6 $T=34040 263840 1 0 $X=33850 $Y=260880
X526 1 2 40 ICV_6 $T=51520 263840 1 0 $X=51330 $Y=260880
X527 1 2 24 ICV_6 $T=51980 220320 0 0 $X=51790 $Y=220080
X528 1 2 42 ICV_6 $T=55660 252960 0 0 $X=55470 $Y=252720
X529 1 2 372 ICV_6 $T=57040 231200 0 0 $X=56850 $Y=230960
X530 1 2 15 ICV_6 $T=57040 236640 0 0 $X=56850 $Y=236400
X531 1 2 26 ICV_6 $T=65320 231200 0 0 $X=65130 $Y=230960
X532 1 2 60 ICV_6 $T=70840 247520 1 0 $X=70650 $Y=244560
X533 1 2 77 ICV_6 $T=97060 263840 1 0 $X=96870 $Y=260880
X534 1 2 414 ICV_6 $T=125580 236640 1 0 $X=125390 $Y=233680
X535 1 2 85 ICV_6 $T=126500 263840 1 0 $X=126310 $Y=260880
X536 1 2 108 ICV_6 $T=135240 252960 0 0 $X=135050 $Y=252720
X537 1 2 422 ICV_6 $T=146280 225760 1 0 $X=146090 $Y=222800
X538 1 2 433 ICV_6 $T=152720 247520 1 0 $X=152530 $Y=244560
X539 1 2 130 ICV_6 $T=167900 247520 0 0 $X=167710 $Y=247280
X540 1 2 445 ICV_6 $T=174800 231200 1 0 $X=174610 $Y=228240
X541 1 2 144 ICV_6 $T=195960 220320 1 0 $X=195770 $Y=217360
X542 1 2 461 ICV_6 $T=203320 231200 1 0 $X=203130 $Y=228240
X543 1 2 123 ICV_6 $T=210220 247520 1 0 $X=210030 $Y=244560
X544 1 2 162 ICV_6 $T=217580 263840 1 0 $X=217390 $Y=260880
X545 1 2 158 ICV_6 $T=238740 236640 0 0 $X=238550 $Y=236400
X546 1 2 495 ICV_6 $T=252540 220320 1 0 $X=252350 $Y=217360
X547 1 2 496 ICV_6 $T=253460 220320 0 0 $X=253270 $Y=220080
X548 1 2 508 ICV_6 $T=276460 247520 0 0 $X=276270 $Y=247280
X549 1 2 516 ICV_6 $T=290260 231200 1 0 $X=290070 $Y=228240
X550 1 2 537 ICV_6 $T=322920 252960 1 0 $X=322730 $Y=250000
X551 1 2 240 ICV_6 $T=323380 220320 1 0 $X=323190 $Y=217360
X552 1 2 536 ICV_6 $T=323840 247520 1 0 $X=323650 $Y=244560
X553 1 2 538 ICV_6 $T=328900 236640 0 0 $X=328710 $Y=236400
X554 1 3 6 ICV_7 $T=7820 220320 1 0 $X=7630 $Y=217360
X555 1 4 350 ICV_7 $T=7820 225760 1 0 $X=7630 $Y=222800
X556 1 3 5 ICV_7 $T=7820 231200 1 0 $X=7630 $Y=228240
X557 1 349 4 ICV_7 $T=7820 236640 0 0 $X=7630 $Y=236400
X558 1 3 4 ICV_7 $T=7820 242080 1 0 $X=7630 $Y=239120
X559 1 3 4 ICV_7 $T=7820 247520 1 0 $X=7630 $Y=244560
X560 1 3 351 ICV_7 $T=7820 252960 1 0 $X=7630 $Y=250000
X561 1 4 352 ICV_7 $T=7820 258400 1 0 $X=7630 $Y=255440
X562 1 7 3 ICV_7 $T=9660 258400 0 0 $X=9470 $Y=258160
X563 1 4 359 ICV_7 $T=20240 247520 0 0 $X=20050 $Y=247280
X564 1 356 360 ICV_7 $T=23460 236640 1 0 $X=23270 $Y=233680
X565 1 19 14 ICV_7 $T=25300 231200 1 0 $X=25110 $Y=228240
X566 1 15 362 ICV_7 $T=26220 236640 0 0 $X=26030 $Y=236400
X567 1 23 24 ICV_7 $T=27600 225760 0 0 $X=27410 $Y=225520
X568 1 363 13 ICV_7 $T=28060 242080 0 0 $X=27870 $Y=241840
X569 1 364 27 ICV_7 $T=29900 236640 0 0 $X=29710 $Y=236400
X570 1 25 22 ICV_7 $T=30360 220320 1 0 $X=30170 $Y=217360
X571 1 27 30 ICV_7 $T=34500 236640 1 0 $X=34310 $Y=233680
X572 1 366 32 ICV_7 $T=38640 231200 1 0 $X=38450 $Y=228240
X573 1 370 14 ICV_7 $T=45080 231200 0 0 $X=44890 $Y=230960
X574 1 19 23 ICV_7 $T=49220 231200 1 0 $X=49030 $Y=228240
X575 1 4 373 ICV_7 $T=51520 242080 0 0 $X=51330 $Y=241840
X576 1 32 369 ICV_7 $T=53360 236640 0 0 $X=53170 $Y=236400
X577 1 4 375 ICV_7 $T=57960 258400 0 0 $X=57770 $Y=258160
X578 1 377 379 ICV_7 $T=63020 220320 0 0 $X=62830 $Y=220080
X579 1 47 380 ICV_7 $T=63940 242080 0 0 $X=63750 $Y=241840
X580 1 48 49 ICV_7 $T=65320 225760 0 0 $X=65130 $Y=225520
X581 1 381 61 ICV_7 $T=67620 236640 0 0 $X=67430 $Y=236400
X582 1 382 65 ICV_7 $T=70380 231200 0 0 $X=70190 $Y=230960
X583 1 61 64 ICV_7 $T=79580 225760 1 0 $X=79390 $Y=222800
X584 1 61 64 ICV_7 $T=80500 231200 0 0 $X=80310 $Y=230960
X585 1 385 389 ICV_7 $T=84180 231200 0 0 $X=83990 $Y=230960
X586 1 393 76 ICV_7 $T=92920 247520 0 0 $X=92730 $Y=247280
X587 1 75 396 ICV_7 $T=92920 252960 0 0 $X=92730 $Y=252720
X588 1 398 400 ICV_7 $T=97980 247520 1 0 $X=97790 $Y=244560
X589 1 79 51 ICV_7 $T=99360 252960 0 0 $X=99170 $Y=252720
X590 1 399 4 ICV_7 $T=99820 225760 0 0 $X=99630 $Y=225520
X591 1 398 401 ICV_7 $T=105340 247520 1 0 $X=105150 $Y=244560
X592 1 402 75 ICV_7 $T=106260 236640 0 0 $X=106070 $Y=236400
X593 1 400 84 ICV_7 $T=107180 247520 0 0 $X=106990 $Y=247280
X594 1 404 398 ICV_7 $T=108560 236640 1 0 $X=108370 $Y=233680
X595 1 405 400 ICV_7 $T=109020 242080 1 0 $X=108830 $Y=239120
X596 1 4 406 ICV_7 $T=111780 252960 0 0 $X=111590 $Y=252720
X597 1 92 85 ICV_7 $T=114080 258400 0 0 $X=113890 $Y=258160
X598 1 93 92 ICV_7 $T=114540 263840 1 0 $X=114350 $Y=260880
X599 1 405 79 ICV_7 $T=120060 242080 1 0 $X=119870 $Y=239120
X600 1 410 4 ICV_7 $T=120060 252960 0 0 $X=119870 $Y=252720
X601 1 75 398 ICV_7 $T=121440 247520 1 0 $X=121250 $Y=244560
X602 1 411 400 ICV_7 $T=121900 231200 0 0 $X=121710 $Y=230960
X603 1 412 94 ICV_7 $T=123280 225760 1 0 $X=123090 $Y=222800
X604 1 4 4 ICV_7 $T=127880 236640 0 0 $X=127690 $Y=236400
X605 1 73 79 ICV_7 $T=132940 231200 0 0 $X=132750 $Y=230960
X606 1 107 112 ICV_7 $T=133860 220320 0 0 $X=133670 $Y=220080
X607 1 109 109 ICV_7 $T=134320 242080 0 0 $X=134130 $Y=241840
X608 1 109 420 ICV_7 $T=140300 252960 0 0 $X=140110 $Y=252720
X609 1 42 115 ICV_7 $T=142140 258400 0 0 $X=141950 $Y=258160
X610 1 428 423 ICV_7 $T=149040 247520 1 0 $X=148850 $Y=244560
X611 1 109 42 ICV_7 $T=149040 252960 0 0 $X=148850 $Y=252720
X612 1 429 431 ICV_7 $T=149500 231200 0 0 $X=149310 $Y=230960
X613 1 428 120 ICV_7 $T=151340 247520 0 0 $X=151150 $Y=247280
X614 1 434 438 ICV_7 $T=154560 236640 0 0 $X=154370 $Y=236400
X615 1 121 123 ICV_7 $T=155480 258400 0 0 $X=155290 $Y=258160
X616 1 437 428 ICV_7 $T=156400 236640 1 0 $X=156210 $Y=233680
X617 1 423 434 ICV_7 $T=156400 242080 1 0 $X=156210 $Y=239120
X618 1 439 440 ICV_7 $T=156400 263840 1 0 $X=156210 $Y=260880
X619 1 425 126 ICV_7 $T=158240 236640 0 0 $X=158050 $Y=236400
X620 1 424 120 ICV_7 $T=160540 247520 0 0 $X=160350 $Y=247280
X621 1 128 434 ICV_7 $T=161460 252960 1 0 $X=161270 $Y=250000
X622 1 119 129 ICV_7 $T=166520 258400 0 0 $X=166330 $Y=258160
X623 1 129 434 ICV_7 $T=169740 252960 0 0 $X=169550 $Y=252720
X624 1 138 448 ICV_7 $T=175260 231200 0 0 $X=175070 $Y=230960
X625 1 450 134 ICV_7 $T=179400 231200 1 0 $X=179210 $Y=228240
X626 1 140 443 ICV_7 $T=179400 236640 1 0 $X=179210 $Y=233680
X627 1 141 142 ICV_7 $T=179400 258400 1 0 $X=179210 $Y=255440
X628 1 451 143 ICV_7 $T=180780 220320 1 0 $X=180590 $Y=217360
X629 1 443 453 ICV_7 $T=182620 236640 0 0 $X=182430 $Y=236400
X630 1 457 147 ICV_7 $T=185380 242080 0 0 $X=185190 $Y=241840
X631 1 146 132 ICV_7 $T=186760 252960 0 0 $X=186570 $Y=252720
X632 1 134 457 ICV_7 $T=190440 236640 0 0 $X=190250 $Y=236400
X633 1 155 352 ICV_7 $T=195500 258400 0 0 $X=195310 $Y=258160
X634 1 4 459 ICV_7 $T=203320 231200 0 0 $X=203130 $Y=230960
X635 1 462 161 ICV_7 $T=204240 236640 0 0 $X=204050 $Y=236400
X636 1 160 164 ICV_7 $T=204700 220320 0 0 $X=204510 $Y=220080
X637 1 463 161 ICV_7 $T=205160 258400 0 0 $X=204970 $Y=258160
X638 1 464 468 ICV_7 $T=205620 252960 0 0 $X=205430 $Y=252720
X639 1 469 469 ICV_7 $T=209300 258400 1 0 $X=209110 $Y=255440
X640 1 467 349 ICV_7 $T=211140 242080 0 0 $X=210950 $Y=241840
X641 1 170 127 ICV_7 $T=212060 263840 1 0 $X=211870 $Y=260880
X642 1 464 172 ICV_7 $T=214820 247520 0 0 $X=214630 $Y=247280
X643 1 473 128 ICV_7 $T=220800 252960 1 0 $X=220610 $Y=250000
X644 1 474 468 ICV_7 $T=220800 258400 0 0 $X=220610 $Y=258160
X645 1 4 476 ICV_7 $T=221260 236640 0 0 $X=221070 $Y=236400
X646 1 468 469 ICV_7 $T=224020 242080 0 0 $X=223830 $Y=241840
X647 1 469 175 ICV_7 $T=224480 258400 0 0 $X=224290 $Y=258160
X648 1 4 477 ICV_7 $T=225860 225760 0 0 $X=225670 $Y=225520
X649 1 478 181 ICV_7 $T=228620 247520 1 0 $X=228430 $Y=244560
X650 1 175 123 ICV_7 $T=232760 258400 1 0 $X=232570 $Y=255440
X651 1 185 483 ICV_7 $T=236440 220320 0 0 $X=236250 $Y=220080
X652 1 488 188 ICV_7 $T=243340 225760 0 0 $X=243150 $Y=225520
X653 1 491 193 ICV_7 $T=245640 231200 1 0 $X=245450 $Y=228240
X654 1 192 487 ICV_7 $T=246560 247520 0 0 $X=246370 $Y=247280
X655 1 486 484 ICV_7 $T=248400 252960 0 0 $X=248210 $Y=252720
X656 1 195 51 ICV_7 $T=248860 220320 1 0 $X=248670 $Y=217360
X657 1 188 193 ICV_7 $T=249780 220320 0 0 $X=249590 $Y=220080
X658 1 190 494 ICV_7 $T=249780 258400 0 0 $X=249590 $Y=258160
X659 1 494 497 ICV_7 $T=252080 252960 0 0 $X=251890 $Y=252720
X660 1 195 195 ICV_7 $T=254380 225760 0 0 $X=254190 $Y=225520
X661 1 501 502 ICV_7 $T=258520 252960 1 0 $X=258330 $Y=250000
X662 1 501 184 ICV_7 $T=258980 258400 1 0 $X=258790 $Y=255440
X663 1 198 481 ICV_7 $T=259900 242080 1 0 $X=259710 $Y=239120
X664 1 486 484 ICV_7 $T=264960 247520 1 0 $X=264770 $Y=244560
X665 1 507 509 ICV_7 $T=268180 231200 0 0 $X=267990 $Y=230960
X666 1 147 512 ICV_7 $T=269560 220320 0 0 $X=269370 $Y=220080
X667 1 512 206 ICV_7 $T=271860 231200 0 0 $X=271670 $Y=230960
X668 1 208 208 ICV_7 $T=275080 225760 0 0 $X=274890 $Y=225520
X669 1 213 216 ICV_7 $T=281060 263840 1 0 $X=280870 $Y=260880
X670 1 512 203 ICV_7 $T=282440 220320 0 0 $X=282250 $Y=220080
X671 1 514 205 ICV_7 $T=283820 236640 1 0 $X=283630 $Y=233680
X672 1 203 512 ICV_7 $T=286580 231200 1 0 $X=286390 $Y=228240
X673 1 206 4 ICV_7 $T=287500 236640 0 0 $X=287310 $Y=236400
X674 1 147 222 ICV_7 $T=287500 258400 0 0 $X=287310 $Y=258160
X675 1 223 179 ICV_7 $T=290720 225760 1 0 $X=290530 $Y=222800
X676 1 192 518 ICV_7 $T=298080 220320 0 0 $X=297890 $Y=220080
X677 1 227 4 ICV_7 $T=302680 225760 0 0 $X=302490 $Y=225520
X678 1 431 522 ICV_7 $T=302680 236640 0 0 $X=302490 $Y=236400
X679 1 230 519 ICV_7 $T=304060 220320 1 0 $X=303870 $Y=217360
X680 1 448 232 ICV_7 $T=305900 258400 0 0 $X=305710 $Y=258160
X681 1 232 521 ICV_7 $T=307280 252960 1 0 $X=307090 $Y=250000
X682 1 521 523 ICV_7 $T=307740 247520 0 0 $X=307550 $Y=247280
X683 1 526 521 ICV_7 $T=310500 236640 0 0 $X=310310 $Y=236400
X684 1 531 239 ICV_7 $T=316020 263840 1 0 $X=315830 $Y=260880
X685 1 532 526 ICV_7 $T=317860 247520 0 0 $X=317670 $Y=247280
X686 1 231 196 ICV_7 $T=319700 220320 1 0 $X=319510 $Y=217360
X687 1 521 521 ICV_7 $T=320160 247520 1 0 $X=319970 $Y=244560
X688 1 431 448 ICV_7 $T=320620 236640 1 0 $X=320430 $Y=233680
X689 1 540 4 ICV_7 $T=326600 231200 0 0 $X=326410 $Y=230960
X690 1 3 4 ICV_7 $T=334880 225760 0 0 $X=334690 $Y=225520
X691 1 3 4 ICV_7 $T=334880 242080 0 0 $X=334690 $Y=241840
X692 1 3 4 ICV_7 $T=335340 220320 0 0 $X=335150 $Y=220080
X693 1 2 3 350 4 2 8 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 220320 0 0 $X=7630 $Y=220080
X694 1 2 3 5 4 2 9 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 231200 0 0 $X=7630 $Y=230960
X695 1 2 3 349 4 2 10 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 242080 0 0 $X=7630 $Y=241840
X696 1 2 3 351 4 2 11 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 247520 0 0 $X=7630 $Y=247280
X697 1 2 3 352 4 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 252960 0 0 $X=7630 $Y=252720
X698 1 2 542 353 4 2 351 1 sky130_fd_sc_hd__dfrtp_4 $T=11500 236640 0 0 $X=11310 $Y=236400
X699 1 2 3 7 4 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=13340 258400 0 0 $X=13150 $Y=258160
X700 1 2 543 354 4 2 21 1 sky130_fd_sc_hd__dfrtp_4 $T=14720 225760 0 0 $X=14530 $Y=225520
X701 1 2 544 359 4 2 20 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 252960 1 0 $X=20970 $Y=250000
X702 1 2 545 365 4 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=33580 258400 1 0 $X=33390 $Y=255440
X703 1 2 546 367 4 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=35880 252960 0 0 $X=35690 $Y=252720
X704 1 2 547 34 4 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=40480 220320 0 0 $X=40290 $Y=220080
X705 1 2 548 373 4 2 47 1 sky130_fd_sc_hd__dfrtp_4 $T=51520 247520 1 0 $X=51330 $Y=244560
X706 1 2 549 375 4 2 55 1 sky130_fd_sc_hd__dfrtp_4 $T=57500 263840 1 0 $X=57310 $Y=260880
X707 1 2 550 376 4 2 63 1 sky130_fd_sc_hd__dfrtp_4 $T=60720 242080 1 0 $X=60530 $Y=239120
X708 1 2 551 378 4 2 60 1 sky130_fd_sc_hd__dfrtp_4 $T=63020 247520 0 0 $X=62830 $Y=247280
X709 1 2 552 67 4 2 71 1 sky130_fd_sc_hd__dfrtp_4 $T=77740 220320 1 0 $X=77550 $Y=217360
X710 1 2 553 386 4 2 70 1 sky130_fd_sc_hd__dfrtp_4 $T=77740 247520 1 0 $X=77550 $Y=244560
X711 1 2 554 390 4 2 77 1 sky130_fd_sc_hd__dfrtp_4 $T=85560 263840 1 0 $X=85370 $Y=260880
X712 1 2 555 392 4 2 74 1 sky130_fd_sc_hd__dfrtp_4 $T=88320 225760 1 0 $X=88130 $Y=222800
X713 1 2 556 72 4 2 80 1 sky130_fd_sc_hd__dfrtp_4 $T=91080 258400 0 0 $X=90890 $Y=258160
X714 1 2 557 394 4 2 81 1 sky130_fd_sc_hd__dfrtp_4 $T=93840 236640 0 0 $X=93650 $Y=236400
X715 1 2 558 399 4 2 90 1 sky130_fd_sc_hd__dfrtp_4 $T=103500 225760 0 0 $X=103310 $Y=225520
X716 1 2 559 406 4 2 100 1 sky130_fd_sc_hd__dfrtp_4 $T=111780 258400 1 0 $X=111590 $Y=255440
X717 1 2 560 407 4 2 97 1 sky130_fd_sc_hd__dfrtp_4 $T=112240 236640 1 0 $X=112050 $Y=233680
X718 1 2 561 412 4 2 106 1 sky130_fd_sc_hd__dfrtp_4 $T=123280 225760 0 0 $X=123090 $Y=225520
X719 1 2 562 413 4 2 108 1 sky130_fd_sc_hd__dfrtp_4 $T=123740 252960 0 0 $X=123550 $Y=252720
X720 1 2 563 415 4 2 113 1 sky130_fd_sc_hd__dfrtp_4 $T=131560 236640 0 0 $X=131370 $Y=236400
X721 1 2 564 416 4 2 114 1 sky130_fd_sc_hd__dfrtp_4 $T=133400 242080 1 0 $X=133210 $Y=239120
X722 1 2 565 417 4 2 116 1 sky130_fd_sc_hd__dfrtp_4 $T=135240 263840 1 0 $X=135050 $Y=260880
X723 1 2 566 422 4 2 6 1 sky130_fd_sc_hd__dfrtp_4 $T=147200 225760 0 0 $X=147010 $Y=225520
X724 1 2 567 432 4 2 124 1 sky130_fd_sc_hd__dfrtp_4 $T=152260 220320 0 0 $X=152070 $Y=220080
X725 1 2 568 436 4 2 130 1 sky130_fd_sc_hd__dfrtp_4 $T=158240 252960 0 0 $X=158050 $Y=252720
X726 1 2 569 133 4 2 135 1 sky130_fd_sc_hd__dfrtp_4 $T=169280 220320 1 0 $X=169090 $Y=217360
X727 1 2 570 447 4 2 352 1 sky130_fd_sc_hd__dfrtp_4 $T=176180 258400 0 0 $X=175990 $Y=258160
X728 1 2 571 452 4 2 149 1 sky130_fd_sc_hd__dfrtp_4 $T=181240 247520 0 0 $X=181050 $Y=247280
X729 1 2 572 459 4 2 167 1 sky130_fd_sc_hd__dfrtp_4 $T=201480 236640 1 0 $X=201290 $Y=233680
X730 1 2 573 461 4 2 166 1 sky130_fd_sc_hd__dfrtp_4 $T=203320 225760 0 0 $X=203130 $Y=225520
X731 1 2 574 460 4 2 349 1 sky130_fd_sc_hd__dfrtp_4 $T=203320 247520 0 0 $X=203130 $Y=247280
X732 1 2 575 476 4 2 181 1 sky130_fd_sc_hd__dfrtp_4 $T=221260 242080 1 0 $X=221070 $Y=239120
X733 1 2 576 477 4 2 183 1 sky130_fd_sc_hd__dfrtp_4 $T=225860 231200 1 0 $X=225670 $Y=228240
X734 1 2 577 479 4 2 187 1 sky130_fd_sc_hd__dfrtp_4 $T=231380 258400 0 0 $X=231190 $Y=258160
X735 1 2 578 482 4 2 191 1 sky130_fd_sc_hd__dfrtp_4 $T=236900 231200 0 0 $X=236710 $Y=230960
X736 1 2 579 491 4 2 194 1 sky130_fd_sc_hd__dfrtp_4 $T=245640 236640 1 0 $X=245450 $Y=233680
X737 1 2 580 489 4 2 189 1 sky130_fd_sc_hd__dfrtp_4 $T=248400 242080 1 0 $X=248210 $Y=239120
X738 1 2 581 510 4 2 211 1 sky130_fd_sc_hd__dfrtp_4 $T=270020 236640 0 0 $X=269830 $Y=236400
X739 1 2 582 506 4 2 210 1 sky130_fd_sc_hd__dfrtp_4 $T=271860 252960 0 0 $X=271670 $Y=252720
X740 1 2 583 505 4 2 214 1 sky130_fd_sc_hd__dfrtp_4 $T=276920 258400 1 0 $X=276730 $Y=255440
X741 1 2 584 221 4 2 225 1 sky130_fd_sc_hd__dfrtp_4 $T=288420 252960 0 0 $X=288230 $Y=252720
X742 1 2 585 517 4 2 226 1 sky130_fd_sc_hd__dfrtp_4 $T=291180 236640 0 0 $X=290990 $Y=236400
X743 1 2 586 529 4 2 235 1 sky130_fd_sc_hd__dfrtp_4 $T=306820 231200 1 0 $X=306630 $Y=228240
X744 1 2 587 520 4 2 238 1 sky130_fd_sc_hd__dfrtp_4 $T=306820 236640 1 0 $X=306630 $Y=233680
X745 1 2 588 234 4 2 350 1 sky130_fd_sc_hd__dfrtp_4 $T=308200 220320 1 0 $X=308010 $Y=217360
X746 1 2 589 537 4 2 541 1 sky130_fd_sc_hd__dfrtp_4 $T=322920 252960 0 0 $X=322730 $Y=252720
X747 1 2 590 535 4 2 244 1 sky130_fd_sc_hd__dfrtp_4 $T=325680 258400 0 0 $X=325490 $Y=258160
X748 1 2 591 540 4 2 243 1 sky130_fd_sc_hd__dfrtp_4 $T=329820 236640 1 0 $X=329630 $Y=233680
X749 1 2 3 242 4 2 249 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 220320 1 0 $X=334690 $Y=217360
X750 1 2 3 246 4 2 250 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 225760 1 0 $X=334690 $Y=222800
X751 1 2 3 247 4 2 251 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 231200 1 0 $X=334690 $Y=228240
X752 1 2 3 541 4 2 252 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 242080 1 0 $X=334690 $Y=239120
X753 1 2 3 248 4 2 253 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 247520 1 0 $X=334690 $Y=244560
X754 1 2 3 245 4 2 254 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 263840 1 0 $X=334690 $Y=260880
X755 1 2 357 ICV_12 $T=21160 236640 1 0 $X=20970 $Y=233680
X756 1 2 356 ICV_12 $T=31280 225760 0 0 $X=31090 $Y=225520
X757 1 2 50 ICV_12 $T=63020 258400 0 0 $X=62830 $Y=258160
X758 1 2 385 ICV_12 $T=77280 225760 1 0 $X=77090 $Y=222800
X759 1 2 68 ICV_12 $T=83260 225760 1 0 $X=83070 $Y=222800
X760 1 2 395 ICV_12 $T=101660 247520 1 0 $X=101470 $Y=244560
X761 1 2 83 ICV_12 $T=112240 263840 1 0 $X=112050 $Y=260880
X762 1 2 98 ICV_12 $T=119140 258400 0 0 $X=118950 $Y=258160
X763 1 2 425 ICV_12 $T=152260 236640 0 0 $X=152070 $Y=236400
X764 1 2 136 ICV_12 $T=180320 220320 0 0 $X=180130 $Y=220080
X765 1 2 171 ICV_12 $T=218500 258400 0 0 $X=218310 $Y=258160
X766 1 2 471 ICV_12 $T=218960 247520 1 0 $X=218770 $Y=244560
X767 1 2 473 ICV_12 $T=227700 242080 0 0 $X=227510 $Y=241840
X768 1 2 479 ICV_12 $T=230460 258400 1 0 $X=230270 $Y=255440
X769 1 2 498 ICV_12 $T=262660 247520 1 0 $X=262470 $Y=244560
X770 1 2 510 ICV_12 $T=270020 236640 1 0 $X=269830 $Y=233680
X771 1 2 117 ICV_12 $T=272780 225760 0 0 $X=272590 $Y=225520
X772 1 2 518 ICV_12 $T=301760 220320 1 0 $X=301570 $Y=217360
X773 1 2 205 ICV_12 $T=301760 220320 0 0 $X=301570 $Y=220080
X774 1 2 156 ICV_12 $T=304980 252960 1 0 $X=304790 $Y=250000
X775 1 2 525 ICV_12 $T=315560 247520 0 0 $X=315370 $Y=247280
X776 1 2 533 ICV_12 $T=317860 247520 1 0 $X=317670 $Y=244560
X777 1 2 238 ICV_12 $T=318320 236640 1 0 $X=318130 $Y=233680
X778 1 2 26 ICV_13 $T=29900 231200 0 0 $X=29710 $Y=230960
X779 1 2 365 ICV_13 $T=31740 252960 1 0 $X=31550 $Y=250000
X780 1 2 26 ICV_13 $T=43240 236640 0 0 $X=43050 $Y=236400
X781 1 2 37 ICV_13 $T=46920 247520 0 0 $X=46730 $Y=247280
X782 1 2 4 ICV_13 $T=73600 242080 0 0 $X=73410 $Y=241840
X783 1 2 4 ICV_13 $T=86020 220320 0 0 $X=85830 $Y=220080
X784 1 2 4 ICV_13 $T=90160 236640 0 0 $X=89970 $Y=236400
X785 1 2 81 ICV_13 $T=99360 242080 0 0 $X=99170 $Y=241840
X786 1 2 46 ICV_13 $T=114080 236640 0 0 $X=113890 $Y=236400
X787 1 2 408 ICV_13 $T=115460 247520 1 0 $X=115270 $Y=244560
X788 1 2 53 ICV_13 $T=126500 247520 0 0 $X=126310 $Y=247280
X789 1 2 416 ICV_13 $T=128340 242080 1 0 $X=128150 $Y=239120
X790 1 2 421 ICV_13 $T=142140 236640 0 0 $X=141950 $Y=236400
X791 1 2 428 ICV_13 $T=147200 236640 1 0 $X=147010 $Y=233680
X792 1 2 431 ICV_13 $T=152260 231200 0 0 $X=152070 $Y=230960
X793 1 2 122 ICV_13 $T=155480 242080 0 0 $X=155290 $Y=241840
X794 1 2 125 ICV_13 $T=156400 258400 1 0 $X=156210 $Y=255440
X795 1 2 442 ICV_13 $T=170200 231200 0 0 $X=170010 $Y=230960
X796 1 2 147 ICV_13 $T=186760 258400 0 0 $X=186570 $Y=258160
X797 1 2 152 ICV_13 $T=189060 225760 0 0 $X=188870 $Y=225520
X798 1 2 4 ICV_13 $T=201480 225760 1 0 $X=201290 $Y=222800
X799 1 2 161 ICV_13 $T=202400 242080 0 0 $X=202210 $Y=241840
X800 1 2 126 ICV_13 $T=229080 263840 1 0 $X=228890 $Y=260880
X801 1 2 492 ICV_13 $T=244720 225760 1 0 $X=244530 $Y=222800
X802 1 2 493 ICV_13 $T=244720 242080 1 0 $X=244530 $Y=239120
X803 1 2 484 ICV_13 $T=251620 247520 1 0 $X=251430 $Y=244560
X804 1 2 4 ICV_13 $T=268180 252960 0 0 $X=267990 $Y=252720
X805 1 2 210 ICV_13 $T=274160 258400 0 0 $X=273970 $Y=258160
X806 1 2 226 ICV_13 $T=292100 242080 0 0 $X=291910 $Y=241840
X807 1 2 534 ICV_13 $T=316940 242080 1 0 $X=316750 $Y=239120
X808 1 2 ICV_14 $T=19780 263840 1 0 $X=19590 $Y=260880
X809 1 2 ICV_14 $T=61640 242080 0 0 $X=61450 $Y=241840
X810 1 2 ICV_14 $T=75900 263840 1 0 $X=75710 $Y=260880
X811 1 2 ICV_14 $T=89700 220320 0 0 $X=89510 $Y=220080
X812 1 2 ICV_14 $T=117760 220320 0 0 $X=117570 $Y=220080
X813 1 2 ICV_14 $T=117760 252960 0 0 $X=117570 $Y=252720
X814 1 2 ICV_14 $T=160080 242080 1 0 $X=159890 $Y=239120
X815 1 2 ICV_14 $T=173880 258400 0 0 $X=173690 $Y=258160
X816 1 2 ICV_14 $T=201940 220320 0 0 $X=201750 $Y=220080
X817 1 2 ICV_14 $T=201940 236640 0 0 $X=201750 $Y=236400
X818 1 2 ICV_14 $T=244260 252960 1 0 $X=244070 $Y=250000
X819 1 2 ICV_14 $T=258060 247520 0 0 $X=257870 $Y=247280
X820 1 2 ICV_14 $T=258060 252960 0 0 $X=257870 $Y=252720
X821 1 2 ICV_14 $T=272320 263840 1 0 $X=272130 $Y=260880
X822 1 2 ICV_14 $T=286120 252960 0 0 $X=285930 $Y=252720
X823 1 2 ICV_14 $T=300380 242080 1 0 $X=300190 $Y=239120
X824 1 13 ICV_15 $T=31740 242080 0 0 $X=31550 $Y=241840
X825 1 4 ICV_15 $T=31740 252960 0 0 $X=31550 $Y=252720
X826 1 4 ICV_15 $T=59800 247520 0 0 $X=59610 $Y=247280
X827 1 68 ICV_15 $T=74060 231200 1 0 $X=73870 $Y=228240
X828 1 384 ICV_15 $T=74060 236640 1 0 $X=73870 $Y=233680
X829 1 391 ICV_15 $T=87860 231200 0 0 $X=87670 $Y=230960
X830 1 82 ICV_15 $T=102120 263840 1 0 $X=101930 $Y=260880
X831 1 400 ICV_15 $T=115920 247520 0 0 $X=115730 $Y=247280
X832 1 106 ICV_15 $T=130180 220320 1 0 $X=129990 $Y=217360
X833 1 415 ICV_15 $T=130180 236640 1 0 $X=129990 $Y=233680
X834 1 79 ICV_15 $T=130180 247520 1 0 $X=129990 $Y=244560
X835 1 409 ICV_15 $T=130180 252960 1 0 $X=129990 $Y=250000
X836 1 4 ICV_15 $T=143980 225760 0 0 $X=143790 $Y=225520
X837 1 434 ICV_15 $T=158240 247520 1 0 $X=158050 $Y=244560
X838 1 436 ICV_15 $T=158240 252960 1 0 $X=158050 $Y=250000
X839 1 135 ICV_15 $T=172040 220320 0 0 $X=171850 $Y=220080
X840 1 144 ICV_15 $T=186300 220320 1 0 $X=186110 $Y=217360
X841 1 145 ICV_15 $T=186300 225760 1 0 $X=186110 $Y=222800
X842 1 453 ICV_15 $T=186300 231200 1 0 $X=186110 $Y=228240
X843 1 4 ICV_15 $T=200100 247520 0 0 $X=199910 $Y=247280
X844 1 179 ICV_15 $T=228160 231200 0 0 $X=227970 $Y=230960
X845 1 4 ICV_15 $T=228160 258400 0 0 $X=227970 $Y=258160
X846 1 511 ICV_15 $T=270480 220320 1 0 $X=270290 $Y=217360
X847 1 515 ICV_15 $T=284280 236640 0 0 $X=284090 $Y=236400
X848 1 218 ICV_15 $T=284280 258400 0 0 $X=284090 $Y=258160
X849 1 141 ICV_15 $T=312340 258400 0 0 $X=312150 $Y=258160
X850 1 2 353 ICV_16 $T=11500 236640 1 0 $X=11310 $Y=233680
X851 1 2 4 ICV_16 $T=12880 263840 1 0 $X=12690 $Y=260880
X852 1 2 4 ICV_16 $T=13340 258400 1 0 $X=13150 $Y=255440
X853 1 2 16 ICV_16 $T=22080 263840 1 0 $X=21890 $Y=260880
X854 1 2 17 ICV_16 $T=23000 220320 1 0 $X=22810 $Y=217360
X855 1 2 20 ICV_16 $T=23920 247520 1 0 $X=23730 $Y=244560
X856 1 2 360 ICV_16 $T=34960 225760 0 0 $X=34770 $Y=225520
X857 1 2 368 ICV_16 $T=37720 247520 1 0 $X=37530 $Y=244560
X858 1 2 369 ICV_16 $T=40020 242080 0 0 $X=39830 $Y=241840
X859 1 2 33 ICV_16 $T=40020 263840 1 0 $X=39830 $Y=260880
X860 1 2 34 ICV_16 $T=40480 220320 1 0 $X=40290 $Y=217360
X861 1 2 370 ICV_16 $T=52900 231200 1 0 $X=52710 $Y=228240
X862 1 2 55 ICV_16 $T=66700 252960 0 0 $X=66510 $Y=252720
X863 1 2 54 ICV_16 $T=70380 258400 0 0 $X=70190 $Y=258160
X864 1 2 69 ICV_16 $T=78200 263840 1 0 $X=78010 $Y=260880
X865 1 2 387 ICV_16 $T=82340 242080 0 0 $X=82150 $Y=241840
X866 1 2 58 ICV_16 $T=92000 231200 1 0 $X=91810 $Y=228240
X867 1 2 74 ICV_16 $T=92460 220320 1 0 $X=92270 $Y=217360
X868 1 2 65 ICV_16 $T=93380 231200 0 0 $X=93190 $Y=230960
X869 1 2 394 ICV_16 $T=93840 236640 1 0 $X=93650 $Y=233680
X870 1 2 397 ICV_16 $T=95220 242080 1 0 $X=95030 $Y=239120
X871 1 2 84 ICV_16 $T=105340 258400 1 0 $X=105150 $Y=255440
X872 1 2 88 ICV_16 $T=109940 220320 1 0 $X=109750 $Y=217360
X873 1 2 96 ICV_16 $T=119140 242080 0 0 $X=118950 $Y=241840
X874 1 2 413 ICV_16 $T=123740 258400 1 0 $X=123550 $Y=255440
X875 1 2 398 ICV_16 $T=125580 231200 1 0 $X=125390 $Y=228240
X876 1 2 100 ICV_16 $T=126500 258400 0 0 $X=126310 $Y=258160
X877 1 2 414 ICV_16 $T=136620 231200 0 0 $X=136430 $Y=230960
X878 1 2 432 ICV_16 $T=152260 220320 1 0 $X=152070 $Y=217360
X879 1 2 6 ICV_16 $T=152260 225760 1 0 $X=152070 $Y=222800
X880 1 2 63 ICV_16 $T=166060 231200 1 0 $X=165870 $Y=228240
X881 1 2 137 ICV_16 $T=177560 252960 0 0 $X=177370 $Y=252720
X882 1 2 452 ICV_16 $T=181240 252960 1 0 $X=181050 $Y=250000
X883 1 2 453 ICV_16 $T=189520 247520 1 0 $X=189330 $Y=244560
X884 1 2 149 ICV_16 $T=192740 247520 0 0 $X=192550 $Y=247280
X885 1 2 89 ICV_16 $T=193660 252960 0 0 $X=193470 $Y=252720
X886 1 2 453 ICV_16 $T=195960 231200 1 0 $X=195770 $Y=228240
X887 1 2 166 ICV_16 $T=213440 220320 0 0 $X=213250 $Y=220080
X888 1 2 167 ICV_16 $T=214820 225760 0 0 $X=214630 $Y=225520
X889 1 2 117 ICV_16 $T=230920 220320 1 0 $X=230730 $Y=217360
X890 1 2 482 ICV_16 $T=236900 236640 1 0 $X=236710 $Y=233680
X891 1 2 4 ICV_16 $T=248400 231200 0 0 $X=248210 $Y=230960
X892 1 2 117 ICV_16 $T=259440 220320 0 0 $X=259250 $Y=220080
X893 1 2 73 ICV_16 $T=260820 225760 1 0 $X=260630 $Y=222800
X894 1 2 182 ICV_16 $T=265880 225760 0 0 $X=265690 $Y=225520
X895 1 2 504 ICV_16 $T=265880 242080 0 0 $X=265690 $Y=241840
X896 1 2 150 ICV_16 $T=287500 225760 0 0 $X=287310 $Y=225520
X897 1 2 517 ICV_16 $T=291640 242080 1 0 $X=291450 $Y=239120
X898 1 2 225 ICV_16 $T=292560 252960 1 0 $X=292370 $Y=250000
X899 1 2 152 ICV_16 $T=293480 220320 1 0 $X=293290 $Y=217360
X900 1 2 516 ICV_16 $T=294860 231200 0 0 $X=294670 $Y=230960
X901 1 2 172 ICV_16 $T=295320 225760 0 0 $X=295130 $Y=225520
X902 1 2 241 ICV_16 $T=320620 225760 1 0 $X=320430 $Y=222800
X903 1 2 539 ICV_16 $T=327520 242080 0 0 $X=327330 $Y=241840
X904 1 2 541 ICV_16 $T=328900 247520 0 0 $X=328710 $Y=247280
X905 1 2 244 ICV_16 $T=334420 252960 0 0 $X=334230 $Y=252720
X906 1 2 245 ICV_16 $T=334880 258400 1 0 $X=334690 $Y=255440
X907 1 2 351 2 356 1 sky130_fd_sc_hd__inv_8 $T=21160 242080 0 0 $X=20970 $Y=241840
X908 1 2 21 2 22 1 sky130_fd_sc_hd__inv_8 $T=23920 225760 1 0 $X=23730 $Y=222800
X909 1 2 20 2 360 1 sky130_fd_sc_hd__inv_8 $T=23920 247520 0 0 $X=23730 $Y=247280
X910 1 2 36 2 366 1 sky130_fd_sc_hd__inv_8 $T=42780 247520 0 0 $X=42590 $Y=247280
X911 1 2 5 2 39 1 sky130_fd_sc_hd__inv_8 $T=49220 220320 1 0 $X=49030 $Y=217360
X912 1 2 37 2 369 1 sky130_fd_sc_hd__inv_8 $T=50600 247520 0 0 $X=50410 $Y=247280
X913 1 2 54 2 56 1 sky130_fd_sc_hd__inv_8 $T=65320 258400 0 0 $X=65130 $Y=258160
X914 1 2 47 2 370 1 sky130_fd_sc_hd__inv_8 $T=65780 247520 1 0 $X=65590 $Y=244560
X915 1 2 55 2 62 1 sky130_fd_sc_hd__inv_8 $T=66700 258400 1 0 $X=66510 $Y=255440
X916 1 2 60 2 382 1 sky130_fd_sc_hd__inv_8 $T=68080 252960 1 0 $X=67890 $Y=250000
X917 1 2 71 2 379 1 sky130_fd_sc_hd__inv_8 $T=81880 220320 0 0 $X=81690 $Y=220080
X918 1 2 70 2 385 1 sky130_fd_sc_hd__inv_8 $T=81880 247520 0 0 $X=81690 $Y=247280
X919 1 2 74 2 389 1 sky130_fd_sc_hd__inv_8 $T=92460 220320 0 0 $X=92270 $Y=220080
X920 1 2 81 2 393 1 sky130_fd_sc_hd__inv_8 $T=103040 242080 0 0 $X=102850 $Y=241840
X921 1 2 80 2 83 1 sky130_fd_sc_hd__inv_8 $T=104420 258400 0 0 $X=104230 $Y=258160
X922 1 2 90 2 94 1 sky130_fd_sc_hd__inv_8 $T=113620 225760 1 0 $X=113430 $Y=222800
X923 1 2 97 2 405 1 sky130_fd_sc_hd__inv_8 $T=119140 231200 1 0 $X=118950 $Y=228240
X924 1 2 100 2 92 1 sky130_fd_sc_hd__inv_8 $T=121440 258400 0 0 $X=121250 $Y=258160
X925 1 2 106 2 111 1 sky130_fd_sc_hd__inv_8 $T=133400 225760 1 0 $X=133210 $Y=222800
X926 1 2 108 2 409 1 sky130_fd_sc_hd__inv_8 $T=133400 258400 1 0 $X=133210 $Y=255440
X927 1 2 112 2 414 1 sky130_fd_sc_hd__inv_8 $T=137540 220320 0 0 $X=137350 $Y=220080
X928 1 2 114 2 423 1 sky130_fd_sc_hd__inv_8 $T=143060 236640 1 0 $X=142870 $Y=233680
X929 1 2 113 2 424 1 sky130_fd_sc_hd__inv_8 $T=147200 236640 0 0 $X=147010 $Y=236400
X930 1 2 6 2 435 1 sky130_fd_sc_hd__inv_8 $T=152260 231200 1 0 $X=152070 $Y=228240
X931 1 2 124 2 442 1 sky130_fd_sc_hd__inv_8 $T=160540 225760 0 0 $X=160350 $Y=225520
X932 1 2 63 2 443 1 sky130_fd_sc_hd__inv_8 $T=166060 231200 0 0 $X=165870 $Y=230960
X933 1 2 130 2 440 1 sky130_fd_sc_hd__inv_8 $T=167900 252960 1 0 $X=167710 $Y=250000
X934 1 2 135 2 449 1 sky130_fd_sc_hd__inv_8 $T=175260 220320 0 0 $X=175070 $Y=220080
X935 1 2 143 2 455 1 sky130_fd_sc_hd__inv_8 $T=182620 220320 0 0 $X=182430 $Y=220080
X936 1 2 149 2 457 1 sky130_fd_sc_hd__inv_8 $T=189520 252960 1 0 $X=189330 $Y=250000
X937 1 2 352 2 155 1 sky130_fd_sc_hd__inv_8 $T=190440 258400 0 0 $X=190250 $Y=258160
X938 1 2 349 2 464 1 sky130_fd_sc_hd__inv_8 $T=206080 242080 0 0 $X=205890 $Y=241840
X939 1 2 166 2 169 1 sky130_fd_sc_hd__inv_8 $T=207920 225760 1 0 $X=207730 $Y=222800
X940 1 2 167 2 466 1 sky130_fd_sc_hd__inv_8 $T=207920 231200 1 0 $X=207730 $Y=228240
X941 1 2 181 2 473 1 sky130_fd_sc_hd__inv_8 $T=231380 242080 0 0 $X=231190 $Y=241840
X942 1 2 183 2 177 1 sky130_fd_sc_hd__inv_8 $T=231840 225760 0 0 $X=231650 $Y=225520
X943 1 2 187 2 487 1 sky130_fd_sc_hd__inv_8 $T=244720 258400 0 0 $X=244530 $Y=258160
X944 1 2 190 2 494 1 sky130_fd_sc_hd__inv_8 $T=245640 263840 1 0 $X=245450 $Y=260880
X945 1 2 194 2 496 1 sky130_fd_sc_hd__inv_8 $T=248400 236640 0 0 $X=248210 $Y=236400
X946 1 2 189 2 498 1 sky130_fd_sc_hd__inv_8 $T=250240 242080 0 0 $X=250050 $Y=241840
X947 1 2 191 2 488 1 sky130_fd_sc_hd__inv_8 $T=259440 231200 0 0 $X=259250 $Y=230960
X948 1 2 211 2 513 1 sky130_fd_sc_hd__inv_8 $T=276460 242080 1 0 $X=276270 $Y=239120
X949 1 2 210 2 501 1 sky130_fd_sc_hd__inv_8 $T=277840 258400 0 0 $X=277650 $Y=258160
X950 1 2 214 2 508 1 sky130_fd_sc_hd__inv_8 $T=281980 252960 1 0 $X=281790 $Y=250000
X951 1 2 225 2 218 1 sky130_fd_sc_hd__inv_8 $T=292560 258400 1 0 $X=292370 $Y=255440
X952 1 2 226 2 516 1 sky130_fd_sc_hd__inv_8 $T=295780 242080 0 0 $X=295590 $Y=241840
X953 1 2 228 2 229 1 sky130_fd_sc_hd__inv_8 $T=301760 263840 1 0 $X=301570 $Y=260880
X954 1 2 235 2 518 1 sky130_fd_sc_hd__inv_8 $T=306360 231200 0 0 $X=306170 $Y=230960
X955 1 2 350 2 237 1 sky130_fd_sc_hd__inv_8 $T=315560 225760 0 0 $X=315370 $Y=225520
X956 1 2 238 2 530 1 sky130_fd_sc_hd__inv_8 $T=315560 236640 0 0 $X=315370 $Y=236400
X957 1 2 541 2 525 1 sky130_fd_sc_hd__inv_8 $T=329820 252960 1 0 $X=329630 $Y=250000
X958 1 2 244 2 532 1 sky130_fd_sc_hd__inv_8 $T=329820 258400 1 0 $X=329630 $Y=255440
X959 1 2 242 2 241 1 sky130_fd_sc_hd__inv_8 $T=330280 220320 0 0 $X=330090 $Y=220080
X960 1 2 243 2 539 1 sky130_fd_sc_hd__inv_8 $T=330280 231200 0 0 $X=330090 $Y=230960
X961 1 2 15 357 2 353 1 sky130_fd_sc_hd__nor2_4 $T=21160 242080 1 0 $X=20970 $Y=239120
X962 1 2 13 363 2 365 1 sky130_fd_sc_hd__nor2_4 $T=32660 247520 1 0 $X=32470 $Y=244560
X963 1 2 13 368 2 367 1 sky130_fd_sc_hd__nor2_4 $T=34960 242080 0 0 $X=34770 $Y=241840
X964 1 2 15 371 2 373 1 sky130_fd_sc_hd__nor2_4 $T=49220 242080 1 0 $X=49030 $Y=239120
X965 1 2 45 374 2 376 1 sky130_fd_sc_hd__nor2_4 $T=60260 252960 1 0 $X=60070 $Y=250000
X966 1 2 15 57 2 59 1 sky130_fd_sc_hd__nor2_4 $T=64860 220320 1 0 $X=64670 $Y=217360
X967 1 2 58 387 2 386 1 sky130_fd_sc_hd__nor2_4 $T=77280 242080 0 0 $X=77090 $Y=241840
X968 1 2 58 388 2 392 1 sky130_fd_sc_hd__nor2_4 $T=91080 225760 0 0 $X=90890 $Y=225520
X969 1 2 75 396 2 390 1 sky130_fd_sc_hd__nor2_4 $T=92920 258400 1 0 $X=92730 $Y=255440
X970 1 2 75 404 2 407 1 sky130_fd_sc_hd__nor2_4 $T=109940 236640 0 0 $X=109750 $Y=236400
X971 1 2 88 110 2 412 1 sky130_fd_sc_hd__nor2_4 $T=133400 220320 1 0 $X=133210 $Y=217360
X972 1 2 109 418 2 416 1 sky130_fd_sc_hd__nor2_4 $T=138000 242080 0 0 $X=137810 $Y=241840
X973 1 2 109 420 2 417 1 sky130_fd_sc_hd__nor2_4 $T=140300 258400 1 0 $X=140110 $Y=255440
X974 1 2 431 429 2 422 1 sky130_fd_sc_hd__nor2_4 $T=151340 236640 1 0 $X=151150 $Y=233680
X975 1 2 431 437 2 432 1 sky130_fd_sc_hd__nor2_4 $T=155940 231200 0 0 $X=155750 $Y=230960
X976 1 2 136 445 2 133 1 sky130_fd_sc_hd__nor2_4 $T=175260 225760 0 0 $X=175070 $Y=225520
X977 1 2 136 451 2 139 1 sky130_fd_sc_hd__nor2_4 $T=178480 225760 1 0 $X=178290 $Y=222800
X978 1 2 141 142 2 447 1 sky130_fd_sc_hd__nor2_4 $T=179400 263840 1 0 $X=179210 $Y=260880
X979 1 2 136 454 2 452 1 sky130_fd_sc_hd__nor2_4 $T=180320 247520 1 0 $X=180130 $Y=244560
X980 1 2 136 151 2 157 1 sky130_fd_sc_hd__nor2_4 $T=190900 220320 1 0 $X=190710 $Y=217360
X981 1 2 161 467 2 460 1 sky130_fd_sc_hd__nor2_4 $T=205160 247520 1 0 $X=204970 $Y=244560
X982 1 2 161 462 2 459 1 sky130_fd_sc_hd__nor2_4 $T=206080 242080 1 0 $X=205890 $Y=239120
X983 1 2 164 160 2 461 1 sky130_fd_sc_hd__nor2_4 $T=208380 220320 0 0 $X=208190 $Y=220080
X984 1 2 136 478 2 479 1 sky130_fd_sc_hd__nor2_4 $T=226320 252960 1 0 $X=226130 $Y=250000
X985 1 2 185 483 2 482 1 sky130_fd_sc_hd__nor2_4 $T=236440 225760 1 0 $X=236250 $Y=222800
X986 1 2 184 480 2 186 1 sky130_fd_sc_hd__nor2_4 $T=236440 258400 1 0 $X=236250 $Y=255440
X987 1 2 206 207 2 204 1 sky130_fd_sc_hd__nor2_4 $T=273700 220320 1 0 $X=273510 $Y=217360
X988 1 2 206 507 2 510 1 sky130_fd_sc_hd__nor2_4 $T=273700 236640 1 0 $X=273510 $Y=233680
X989 1 2 206 515 2 517 1 sky130_fd_sc_hd__nor2_4 $T=286580 242080 1 0 $X=286390 $Y=239120
X990 1 2 431 522 2 520 1 sky130_fd_sc_hd__nor2_4 $T=302680 242080 1 0 $X=302490 $Y=239120
X991 1 2 227 524 2 529 1 sky130_fd_sc_hd__nor2_4 $T=306360 225760 0 0 $X=306170 $Y=225520
X992 1 2 227 236 2 234 1 sky130_fd_sc_hd__nor2_4 $T=310960 225760 1 0 $X=310770 $Y=222800
X993 1 2 431 533 2 535 1 sky130_fd_sc_hd__nor2_4 $T=315560 252960 0 0 $X=315370 $Y=252720
X994 1 2 141 531 2 537 1 sky130_fd_sc_hd__nor2_4 $T=315560 258400 0 0 $X=315370 $Y=258160
X995 1 2 431 538 2 540 1 sky130_fd_sc_hd__nor2_4 $T=320620 242080 1 0 $X=320430 $Y=239120
X996 1 2 356 19 14 355 2 357 1 sky130_fd_sc_hd__o22a_4 $T=23460 231200 0 0 $X=23270 $Y=230960
X997 1 2 360 19 14 358 2 361 1 sky130_fd_sc_hd__o22a_4 $T=27140 236640 1 0 $X=26950 $Y=233680
X998 1 2 366 27 30 364 2 363 1 sky130_fd_sc_hd__o22a_4 $T=36340 242080 1 0 $X=36150 $Y=239120
X999 1 2 369 27 30 362 2 368 1 sky130_fd_sc_hd__o22a_4 $T=36800 236640 0 0 $X=36610 $Y=236400
X1000 1 2 370 19 14 372 2 371 1 sky130_fd_sc_hd__o22a_4 $T=49220 236640 1 0 $X=49030 $Y=233680
X1001 1 2 379 64 61 377 2 383 1 sky130_fd_sc_hd__o22a_4 $T=71300 220320 0 0 $X=71110 $Y=220080
X1002 1 2 382 64 61 381 2 380 1 sky130_fd_sc_hd__o22a_4 $T=71300 236640 0 0 $X=71110 $Y=236400
X1003 1 2 385 64 61 384 2 387 1 sky130_fd_sc_hd__o22a_4 $T=77280 236640 1 0 $X=77090 $Y=233680
X1004 1 2 389 64 61 391 2 388 1 sky130_fd_sc_hd__o22a_4 $T=79580 225760 0 0 $X=79390 $Y=225520
X1005 1 2 393 398 400 395 2 397 1 sky130_fd_sc_hd__o22a_4 $T=99820 247520 0 0 $X=99630 $Y=247280
X1006 1 2 84 398 400 401 2 396 1 sky130_fd_sc_hd__o22a_4 $T=105340 252960 1 0 $X=105150 $Y=250000
X1007 1 2 405 398 400 402 2 404 1 sky130_fd_sc_hd__o22a_4 $T=112700 242080 1 0 $X=112510 $Y=239120
X1008 1 2 94 102 104 101 2 403 1 sky130_fd_sc_hd__o22a_4 $T=120060 220320 1 0 $X=119870 $Y=217360
X1009 1 2 409 398 400 410 2 408 1 sky130_fd_sc_hd__o22a_4 $T=120060 247520 0 0 $X=119870 $Y=247280
X1010 1 2 414 398 400 411 2 105 1 sky130_fd_sc_hd__o22a_4 $T=125580 231200 0 0 $X=125390 $Y=230960
X1011 1 2 119 117 115 426 2 118 1 sky130_fd_sc_hd__o22a_4 $T=147200 258400 0 0 $X=147010 $Y=258160
X1012 1 2 424 428 425 421 2 419 1 sky130_fd_sc_hd__o22a_4 $T=149040 242080 1 0 $X=148850 $Y=239120
X1013 1 2 423 428 425 433 2 418 1 sky130_fd_sc_hd__o22a_4 $T=149040 242080 0 0 $X=148850 $Y=241840
X1014 1 2 120 428 425 427 2 420 1 sky130_fd_sc_hd__o22a_4 $T=149500 252960 1 0 $X=149310 $Y=250000
X1015 1 2 440 125 121 439 2 430 1 sky130_fd_sc_hd__o22a_4 $T=159160 258400 0 0 $X=158970 $Y=258160
X1016 1 2 435 428 425 441 2 429 1 sky130_fd_sc_hd__o22a_4 $T=161460 236640 1 0 $X=161270 $Y=233680
X1017 1 2 442 428 425 438 2 437 1 sky130_fd_sc_hd__o22a_4 $T=161920 236640 0 0 $X=161730 $Y=236400
X1018 1 2 443 134 446 444 2 374 1 sky130_fd_sc_hd__o22a_4 $T=175260 236640 0 0 $X=175070 $Y=236400
X1019 1 2 449 134 446 456 2 445 1 sky130_fd_sc_hd__o22a_4 $T=181240 231200 0 0 $X=181050 $Y=230960
X1020 1 2 455 134 446 450 2 451 1 sky130_fd_sc_hd__o22a_4 $T=182620 225760 0 0 $X=182430 $Y=225520
X1021 1 2 144 134 446 154 2 151 1 sky130_fd_sc_hd__o22a_4 $T=189520 225760 1 0 $X=189330 $Y=222800
X1022 1 2 457 134 446 458 2 454 1 sky130_fd_sc_hd__o22a_4 $T=189520 242080 1 0 $X=189330 $Y=239120
X1023 1 2 464 469 468 465 2 467 1 sky130_fd_sc_hd__o22a_4 $T=209300 252960 0 0 $X=209110 $Y=252720
X1024 1 2 466 469 468 470 2 462 1 sky130_fd_sc_hd__o22a_4 $T=210220 236640 0 0 $X=210030 $Y=236400
X1025 1 2 170 469 468 171 2 463 1 sky130_fd_sc_hd__o22a_4 $T=211140 258400 0 0 $X=210950 $Y=258160
X1026 1 2 473 469 468 472 2 471 1 sky130_fd_sc_hd__o22a_4 $T=221260 247520 1 0 $X=221070 $Y=244560
X1027 1 2 175 469 468 474 2 173 1 sky130_fd_sc_hd__o22a_4 $T=222640 263840 1 0 $X=222450 $Y=260880
X1028 1 2 177 176 180 174 2 475 1 sky130_fd_sc_hd__o22a_4 $T=223560 220320 1 0 $X=223370 $Y=217360
X1029 1 2 487 484 486 485 2 478 1 sky130_fd_sc_hd__o22a_4 $T=241040 252960 0 0 $X=240850 $Y=252720
X1030 1 2 488 193 188 492 2 483 1 sky130_fd_sc_hd__o22a_4 $T=247020 225760 0 0 $X=246830 $Y=225520
X1031 1 2 494 484 486 497 2 480 1 sky130_fd_sc_hd__o22a_4 $T=247940 258400 1 0 $X=247750 $Y=255440
X1032 1 2 496 193 188 495 2 490 1 sky130_fd_sc_hd__o22a_4 $T=248400 225760 1 0 $X=248210 $Y=222800
X1033 1 2 498 484 486 500 2 493 1 sky130_fd_sc_hd__o22a_4 $T=255300 247520 1 0 $X=255110 $Y=244560
X1034 1 2 501 484 486 499 2 503 1 sky130_fd_sc_hd__o22a_4 $T=262200 252960 1 0 $X=262010 $Y=250000
X1035 1 2 508 484 486 504 2 502 1 sky130_fd_sc_hd__o22a_4 $T=264960 247520 0 0 $X=264770 $Y=247280
X1036 1 2 208 512 203 511 2 207 1 sky130_fd_sc_hd__o22a_4 $T=275080 220320 0 0 $X=274890 $Y=220080
X1037 1 2 513 512 203 509 2 507 1 sky130_fd_sc_hd__o22a_4 $T=276000 231200 0 0 $X=275810 $Y=230960
X1038 1 2 217 512 203 219 2 215 1 sky130_fd_sc_hd__o22a_4 $T=281980 220320 1 0 $X=281790 $Y=217360
X1039 1 2 223 512 203 224 2 220 1 sky130_fd_sc_hd__o22a_4 $T=287500 220320 0 0 $X=287310 $Y=220080
X1040 1 2 516 512 203 514 2 515 1 sky130_fd_sc_hd__o22a_4 $T=287500 231200 0 0 $X=287310 $Y=230960
X1041 1 2 518 231 230 519 2 524 1 sky130_fd_sc_hd__o22a_4 $T=304060 220320 0 0 $X=303870 $Y=220080
X1042 1 2 232 521 526 528 2 233 1 sky130_fd_sc_hd__o22a_4 $T=309120 258400 1 0 $X=308930 $Y=255440
X1043 1 2 530 521 526 527 2 522 1 sky130_fd_sc_hd__o22a_4 $T=310500 242080 1 0 $X=310310 $Y=239120
X1044 1 2 525 521 526 523 2 531 1 sky130_fd_sc_hd__o22a_4 $T=311420 252960 1 0 $X=311230 $Y=250000
X1045 1 2 539 521 526 534 2 538 1 sky130_fd_sc_hd__o22a_4 $T=320160 242080 0 0 $X=319970 $Y=241840
X1046 1 2 532 521 526 536 2 533 1 sky130_fd_sc_hd__o22a_4 $T=321540 247520 0 0 $X=321350 $Y=247280
X1047 1 2 24 2 38 1 sky130_fd_sc_hd__buf_1 $T=49220 225760 1 0 $X=49030 $Y=222800
X1048 1 2 35 2 44 1 sky130_fd_sc_hd__buf_1 $T=55660 225760 0 0 $X=55470 $Y=225520
X1049 1 2 42 2 45 1 sky130_fd_sc_hd__buf_1 $T=55660 258400 1 0 $X=55470 $Y=255440
X1050 1 2 43 2 46 1 sky130_fd_sc_hd__buf_1 $T=56580 220320 0 0 $X=56390 $Y=220080
X1051 1 2 48 2 51 1 sky130_fd_sc_hd__buf_1 $T=63020 225760 0 0 $X=62830 $Y=225520
X1052 1 2 26 2 52 1 sky130_fd_sc_hd__buf_1 $T=63020 231200 0 0 $X=62830 $Y=230960
X1053 1 2 49 2 53 1 sky130_fd_sc_hd__buf_1 $T=63480 231200 1 0 $X=63290 $Y=228240
X1054 1 2 65 2 73 1 sky130_fd_sc_hd__buf_1 $T=91080 231200 0 0 $X=90890 $Y=230960
X1055 1 2 89 2 79 1 sky130_fd_sc_hd__buf_1 $T=112700 231200 1 0 $X=112510 $Y=228240
X1056 1 2 91 2 398 1 sky130_fd_sc_hd__buf_1 $T=114080 247520 1 0 $X=113890 $Y=244560
X1057 1 2 96 2 400 1 sky130_fd_sc_hd__buf_1 $T=119140 247520 1 0 $X=118950 $Y=244560
X1058 1 2 107 2 75 1 sky130_fd_sc_hd__buf_1 $T=131560 220320 0 0 $X=131370 $Y=220080
X1059 1 2 42 2 109 1 sky130_fd_sc_hd__buf_1 $T=139840 258400 0 0 $X=139650 $Y=258160
X1060 1 2 117 2 102 1 sky130_fd_sc_hd__buf_1 $T=147200 220320 1 0 $X=147010 $Y=217360
X1061 1 2 42 2 431 1 sky130_fd_sc_hd__buf_1 $T=152720 252960 0 0 $X=152530 $Y=252720
X1062 1 2 131 2 428 1 sky130_fd_sc_hd__buf_1 $T=168820 242080 0 0 $X=168630 $Y=241840
X1063 1 2 132 2 434 1 sky130_fd_sc_hd__buf_1 $T=169740 263840 1 0 $X=169550 $Y=260880
X1064 1 2 137 2 425 1 sky130_fd_sc_hd__buf_1 $T=175260 242080 0 0 $X=175070 $Y=241840
X1065 1 2 137 2 121 1 sky130_fd_sc_hd__buf_1 $T=175260 252960 0 0 $X=175070 $Y=252720
X1066 1 2 131 2 125 1 sky130_fd_sc_hd__buf_1 $T=175720 252960 1 0 $X=175530 $Y=250000
X1067 1 2 132 2 448 1 sky130_fd_sc_hd__buf_1 $T=189520 258400 1 0 $X=189330 $Y=255440
X1068 1 2 146 2 453 1 sky130_fd_sc_hd__buf_1 $T=190440 252960 0 0 $X=190250 $Y=252720
X1069 1 2 153 2 446 1 sky130_fd_sc_hd__buf_1 $T=191360 231200 0 0 $X=191170 $Y=230960
X1070 1 2 89 2 123 1 sky130_fd_sc_hd__buf_1 $T=193660 258400 1 0 $X=193470 $Y=255440
X1071 1 2 158 2 134 1 sky130_fd_sc_hd__buf_1 $T=196420 231200 0 0 $X=196230 $Y=230960
X1072 1 2 89 2 159 1 sky130_fd_sc_hd__buf_1 $T=201940 220320 1 0 $X=201750 $Y=217360
X1073 1 2 172 2 161 1 sky130_fd_sc_hd__buf_1 $T=217580 252960 1 0 $X=217390 $Y=250000
X1074 1 2 117 2 176 1 sky130_fd_sc_hd__buf_1 $T=231380 220320 0 0 $X=231190 $Y=220080
X1075 1 2 179 2 468 1 sky130_fd_sc_hd__buf_1 $T=231380 231200 0 0 $X=231190 $Y=230960
X1076 1 2 182 2 469 1 sky130_fd_sc_hd__buf_1 $T=231840 236640 1 0 $X=231650 $Y=233680
X1077 1 2 146 2 481 1 sky130_fd_sc_hd__buf_1 $T=235980 252960 0 0 $X=235790 $Y=252720
X1078 1 2 158 2 484 1 sky130_fd_sc_hd__buf_1 $T=238740 242080 1 0 $X=238550 $Y=239120
X1079 1 2 153 2 486 1 sky130_fd_sc_hd__buf_1 $T=244260 242080 0 0 $X=244070 $Y=241840
X1080 1 2 117 2 193 1 sky130_fd_sc_hd__buf_1 $T=258520 225760 1 0 $X=258330 $Y=222800
X1081 1 2 182 2 117 1 sky130_fd_sc_hd__buf_1 $T=261740 231200 1 0 $X=261550 $Y=228240
X1082 1 2 117 2 512 1 sky130_fd_sc_hd__buf_1 $T=273700 231200 1 0 $X=273510 $Y=228240
X1083 1 2 172 2 206 1 sky130_fd_sc_hd__buf_1 $T=281520 236640 1 0 $X=281330 $Y=233680
X1084 1 2 179 2 203 1 sky130_fd_sc_hd__buf_1 $T=288420 225760 1 0 $X=288230 $Y=222800
X1085 1 2 172 2 227 1 sky130_fd_sc_hd__buf_1 $T=295320 231200 1 0 $X=295130 $Y=228240
X1086 1 2 131 2 521 1 sky130_fd_sc_hd__buf_1 $T=302220 247520 0 0 $X=302030 $Y=247280
X1087 1 2 137 2 526 1 sky130_fd_sc_hd__buf_1 $T=305440 247520 1 0 $X=305250 $Y=244560
X1088 1 2 24 356 23 2 355 1 sky130_fd_sc_hd__o21a_4 $T=29440 231200 1 0 $X=29250 $Y=228240
X1089 1 2 31 22 32 2 28 1 sky130_fd_sc_hd__o21a_4 $T=34040 220320 1 0 $X=33850 $Y=217360
X1090 1 2 26 360 23 2 358 1 sky130_fd_sc_hd__o21a_4 $T=34960 231200 0 0 $X=34770 $Y=230960
X1091 1 2 35 366 32 2 364 1 sky130_fd_sc_hd__o21a_4 $T=38640 236640 1 0 $X=38450 $Y=233680
X1092 1 2 26 369 32 2 362 1 sky130_fd_sc_hd__o21a_4 $T=46920 236640 0 0 $X=46730 $Y=236400
X1093 1 2 35 370 23 2 372 1 sky130_fd_sc_hd__o21a_4 $T=50600 231200 0 0 $X=50410 $Y=230960
X1094 1 2 43 379 23 2 377 1 sky130_fd_sc_hd__o21a_4 $T=66700 225760 1 0 $X=66510 $Y=222800
X1095 1 2 65 382 68 2 381 1 sky130_fd_sc_hd__o21a_4 $T=74060 231200 0 0 $X=73870 $Y=230960
X1096 1 2 48 385 68 2 384 1 sky130_fd_sc_hd__o21a_4 $T=77280 231200 1 0 $X=77090 $Y=228240
X1097 1 2 49 389 68 2 391 1 sky130_fd_sc_hd__o21a_4 $T=85560 231200 1 0 $X=85370 $Y=228240
X1098 1 2 76 393 78 2 395 1 sky130_fd_sc_hd__o21a_4 $T=94760 252960 1 0 $X=94570 $Y=250000
X1099 1 2 51 84 79 2 401 1 sky130_fd_sc_hd__o21a_4 $T=103040 252960 0 0 $X=102850 $Y=252720
X1100 1 2 98 92 85 2 95 1 sky130_fd_sc_hd__o21a_4 $T=118680 263840 1 0 $X=118490 $Y=260880
X1101 1 2 46 405 79 2 402 1 sky130_fd_sc_hd__o21a_4 $T=119140 236640 0 0 $X=118950 $Y=236400
X1102 1 2 103 94 99 2 101 1 sky130_fd_sc_hd__o21a_4 $T=122360 220320 0 0 $X=122170 $Y=220080
X1103 1 2 53 409 79 2 410 1 sky130_fd_sc_hd__o21a_4 $T=130180 247520 0 0 $X=129990 $Y=247280
X1104 1 2 73 414 79 2 411 1 sky130_fd_sc_hd__o21a_4 $T=133400 236640 1 0 $X=133210 $Y=233680
X1105 1 2 127 423 434 2 433 1 sky130_fd_sc_hd__o21a_4 $T=159160 242080 0 0 $X=158970 $Y=241840
X1106 1 2 122 424 434 2 421 1 sky130_fd_sc_hd__o21a_4 $T=161460 247520 1 0 $X=161270 $Y=244560
X1107 1 2 128 120 434 2 427 1 sky130_fd_sc_hd__o21a_4 $T=161460 258400 1 0 $X=161270 $Y=255440
X1108 1 2 129 119 123 2 426 1 sky130_fd_sc_hd__o21a_4 $T=161460 263840 1 0 $X=161270 $Y=260880
X1109 1 2 126 435 434 2 441 1 sky130_fd_sc_hd__o21a_4 $T=162380 242080 1 0 $X=162190 $Y=239120
X1110 1 2 129 440 434 2 439 1 sky130_fd_sc_hd__o21a_4 $T=169740 258400 1 0 $X=169550 $Y=255440
X1111 1 2 138 442 448 2 438 1 sky130_fd_sc_hd__o21a_4 $T=172960 236640 1 0 $X=172770 $Y=233680
X1112 1 2 140 443 453 2 444 1 sky130_fd_sc_hd__o21a_4 $T=178020 242080 1 0 $X=177830 $Y=239120
X1113 1 2 147 457 453 2 458 1 sky130_fd_sc_hd__o21a_4 $T=189060 242080 0 0 $X=188870 $Y=241840
X1114 1 2 145 449 453 2 456 1 sky130_fd_sc_hd__o21a_4 $T=189520 231200 1 0 $X=189330 $Y=228240
X1115 1 2 147 155 156 2 148 1 sky130_fd_sc_hd__o21a_4 $T=189520 263840 1 0 $X=189330 $Y=260880
X1116 1 2 150 144 453 2 154 1 sky130_fd_sc_hd__o21a_4 $T=191820 220320 0 0 $X=191630 $Y=220080
X1117 1 2 152 455 453 2 450 1 sky130_fd_sc_hd__o21a_4 $T=192740 225760 0 0 $X=192550 $Y=225520
X1118 1 2 168 169 99 2 163 1 sky130_fd_sc_hd__o21a_4 $T=207000 220320 1 0 $X=206810 $Y=217360
X1119 1 2 122 464 123 2 465 1 sky130_fd_sc_hd__o21a_4 $T=207000 252960 1 0 $X=206810 $Y=250000
X1120 1 2 138 466 159 2 470 1 sky130_fd_sc_hd__o21a_4 $T=211140 231200 0 0 $X=210950 $Y=230960
X1121 1 2 128 473 123 2 472 1 sky130_fd_sc_hd__o21a_4 $T=220800 247520 0 0 $X=220610 $Y=247280
X1122 1 2 52 177 178 2 174 1 sky130_fd_sc_hd__o21a_4 $T=226320 225760 1 0 $X=226130 $Y=222800
X1123 1 2 126 175 123 2 474 1 sky130_fd_sc_hd__o21a_4 $T=232760 263840 1 0 $X=232570 $Y=260880
X1124 1 2 192 487 481 2 485 1 sky130_fd_sc_hd__o21a_4 $T=246560 252960 1 0 $X=246370 $Y=250000
X1125 1 2 53 496 195 2 495 1 sky130_fd_sc_hd__o21a_4 $T=251620 231200 1 0 $X=251430 $Y=228240
X1126 1 2 196 494 481 2 497 1 sky130_fd_sc_hd__o21a_4 $T=253460 263840 1 0 $X=253270 $Y=260880
X1127 1 2 46 200 195 2 197 1 sky130_fd_sc_hd__o21a_4 $T=258520 220320 1 0 $X=258330 $Y=217360
X1128 1 2 73 488 195 2 492 1 sky130_fd_sc_hd__o21a_4 $T=259440 225760 0 0 $X=259250 $Y=225520
X1129 1 2 198 498 481 2 500 1 sky130_fd_sc_hd__o21a_4 $T=259440 242080 0 0 $X=259250 $Y=241840
X1130 1 2 199 501 481 2 499 1 sky130_fd_sc_hd__o21a_4 $T=262660 252960 0 0 $X=262470 $Y=252720
X1131 1 2 202 508 481 2 504 1 sky130_fd_sc_hd__o21a_4 $T=273700 252960 1 0 $X=273510 $Y=250000
X1132 1 2 147 208 205 2 511 1 sky130_fd_sc_hd__o21a_4 $T=276000 225760 1 0 $X=275810 $Y=222800
X1133 1 2 145 513 205 2 509 1 sky130_fd_sc_hd__o21a_4 $T=279220 231200 1 0 $X=279030 $Y=228240
X1134 1 2 147 218 222 2 213 1 sky130_fd_sc_hd__o21a_4 $T=285200 263840 1 0 $X=285010 $Y=260880
X1135 1 2 150 516 205 2 514 1 sky130_fd_sc_hd__o21a_4 $T=287500 236640 1 0 $X=287310 $Y=233680
X1136 1 2 192 518 205 2 519 1 sky130_fd_sc_hd__o21a_4 $T=301760 225760 1 0 $X=301570 $Y=222800
X1137 1 2 192 525 156 2 523 1 sky130_fd_sc_hd__o21a_4 $T=304980 252960 0 0 $X=304790 $Y=252720
X1138 1 2 198 232 448 2 528 1 sky130_fd_sc_hd__o21a_4 $T=309580 263840 1 0 $X=309390 $Y=260880
X1139 1 2 196 530 448 2 527 1 sky130_fd_sc_hd__o21a_4 $T=311420 247520 1 0 $X=311230 $Y=244560
X1140 1 2 202 532 448 2 536 1 sky130_fd_sc_hd__o21a_4 $T=319240 258400 1 0 $X=319050 $Y=255440
X1141 1 2 196 241 159 2 240 1 sky130_fd_sc_hd__o21a_4 $T=320620 220320 0 0 $X=320430 $Y=220080
X1142 1 2 199 539 448 2 534 1 sky130_fd_sc_hd__o21a_4 $T=322460 236640 0 0 $X=322270 $Y=236400
X1143 1 2 355 14 ICV_21 $T=18400 231200 0 0 $X=18210 $Y=230960
X1144 1 2 358 19 ICV_21 $T=20240 231200 1 0 $X=20050 $Y=228240
X1145 1 2 4 367 ICV_21 $T=34500 252960 1 0 $X=34310 $Y=250000
X1146 1 2 374 45 ICV_21 $T=54740 247520 0 0 $X=54550 $Y=247280
X1147 1 2 386 58 ICV_21 $T=76360 242080 1 0 $X=76170 $Y=239120
X1148 1 2 390 4 ICV_21 $T=82340 258400 0 0 $X=82150 $Y=258160
X1149 1 2 4 407 ICV_21 $T=110860 231200 0 0 $X=110670 $Y=230960
X1150 1 2 113 424 ICV_21 $T=143980 242080 1 0 $X=143790 $Y=239120
X1151 1 2 426 117 ICV_21 $T=145820 263840 1 0 $X=145630 $Y=260880
X1152 1 2 427 425 ICV_21 $T=146280 247520 0 0 $X=146090 $Y=247280
X1153 1 2 444 446 ICV_21 $T=171580 242080 1 0 $X=171390 $Y=239120
X1154 1 2 458 446 ICV_21 $T=185380 236640 0 0 $X=185190 $Y=236400
X1155 1 2 446 150 ICV_21 $T=186760 220320 0 0 $X=186570 $Y=220080
X1156 1 2 466 159 ICV_21 $T=206080 231200 0 0 $X=205890 $Y=230960
X1157 1 2 489 4 ICV_21 $T=243340 236640 0 0 $X=243150 $Y=236400
X1158 1 2 202 481 ICV_21 $T=271400 247520 0 0 $X=271210 $Y=247280
X1159 1 2 205 513 ICV_21 $T=277840 225760 0 0 $X=277650 $Y=225520
X1160 1 2 205 223 ICV_21 $T=288420 220320 1 0 $X=288230 $Y=217360
X1161 1 2 520 4 ICV_21 $T=301300 231200 0 0 $X=301110 $Y=230960
X1162 1 2 527 530 ICV_21 $T=305440 236640 0 0 $X=305250 $Y=236400
X1163 1 2 202 448 ICV_21 $T=317860 252960 1 0 $X=317670 $Y=250000
X1164 1 2 3 4 ICV_21 $T=333500 236640 0 0 $X=333310 $Y=236400
X1165 1 2 36 ICV_22 $T=39560 247520 0 0 $X=39370 $Y=247280
X1166 1 2 4 ICV_22 $T=86480 258400 0 0 $X=86290 $Y=258160
X1167 1 2 91 ICV_22 $T=112700 242080 0 0 $X=112510 $Y=241840
X1168 1 2 4 ICV_22 $T=120060 225760 0 0 $X=119870 $Y=225520
X1169 1 2 131 ICV_22 $T=174340 247520 0 0 $X=174150 $Y=247280
X1170 1 2 446 ICV_22 $T=178020 231200 0 0 $X=177830 $Y=230960
X1171 1 2 446 ICV_22 $T=179400 225760 0 0 $X=179210 $Y=225520
X1172 1 2 468 ICV_22 $T=207000 236640 0 0 $X=206810 $Y=236400
X1173 1 2 468 ICV_22 $T=207920 258400 0 0 $X=207730 $Y=258160
X1174 1 2 123 ICV_22 $T=217580 247520 0 0 $X=217390 $Y=247280
X1175 1 2 52 ICV_22 $T=223100 225760 1 0 $X=222910 $Y=222800
X1176 1 2 484 ICV_22 $T=239660 247520 0 0 $X=239470 $Y=247280
X1177 1 2 153 ICV_22 $T=241040 242080 0 0 $X=240850 $Y=241840
X1178 1 2 53 ICV_22 $T=248400 231200 1 0 $X=248210 $Y=228240
X1179 1 2 191 ICV_22 $T=254840 231200 0 0 $X=254650 $Y=230960
X1180 1 2 205 ICV_22 $T=272780 225760 1 0 $X=272590 $Y=222800
X1181 1 2 212 ICV_22 $T=276000 263840 1 0 $X=275810 $Y=260880
X1182 1 2 512 ICV_22 $T=285200 225760 1 0 $X=285010 $Y=222800
X1183 1 2 228 ICV_22 $T=299460 258400 0 0 $X=299270 $Y=258160
X1184 1 2 528 ICV_22 $T=305900 258400 1 0 $X=305710 $Y=255440
X1185 1 2 4 ICV_22 $T=319700 252960 0 0 $X=319510 $Y=252720
X1186 1 2 243 ICV_22 $T=328900 231200 1 0 $X=328710 $Y=228240
X1187 1 2 ICV_23 $T=18400 252960 0 0 $X=18210 $Y=252720
X1188 1 2 ICV_23 $T=20240 258400 1 0 $X=20050 $Y=255440
X1189 1 2 ICV_23 $T=28060 225760 1 0 $X=27870 $Y=222800
X1190 1 2 ICV_23 $T=34040 258400 0 0 $X=33850 $Y=258160
X1191 1 2 ICV_23 $T=41400 225760 0 0 $X=41210 $Y=225520
X1192 1 2 ICV_23 $T=48300 252960 1 0 $X=48110 $Y=250000
X1193 1 2 ICV_23 $T=50600 225760 1 0 $X=50410 $Y=222800
X1194 1 2 ICV_23 $T=53360 220320 1 0 $X=53170 $Y=217360
X1195 1 2 ICV_23 $T=55660 236640 1 0 $X=55470 $Y=233680
X1196 1 2 ICV_23 $T=73140 252960 0 0 $X=72950 $Y=252720
X1197 1 2 ICV_23 $T=76360 252960 1 0 $X=76170 $Y=250000
X1198 1 2 ICV_23 $T=76360 258400 1 0 $X=76170 $Y=255440
X1199 1 2 ICV_23 $T=77740 236640 0 0 $X=77550 $Y=236400
X1200 1 2 ICV_23 $T=80500 242080 1 0 $X=80310 $Y=239120
X1201 1 2 ICV_23 $T=96600 220320 0 0 $X=96410 $Y=220080
X1202 1 2 ICV_23 $T=99820 231200 0 0 $X=99630 $Y=230960
X1203 1 2 ICV_23 $T=132480 231200 1 0 $X=132290 $Y=228240
X1204 1 2 ICV_23 $T=132480 252960 1 0 $X=132290 $Y=250000
X1205 1 2 ICV_23 $T=160540 225760 1 0 $X=160350 $Y=222800
X1206 1 2 ICV_23 $T=166980 247520 1 0 $X=166790 $Y=244560
X1207 1 2 ICV_23 $T=188600 236640 1 0 $X=188410 $Y=233680
X1208 1 2 ICV_23 $T=193660 252960 1 0 $X=193470 $Y=250000
X1209 1 2 ICV_23 $T=195040 258400 1 0 $X=194850 $Y=255440
X1210 1 2 ICV_23 $T=215740 252960 0 0 $X=215550 $Y=252720
X1211 1 2 ICV_23 $T=216660 231200 0 0 $X=216470 $Y=230960
X1212 1 2 ICV_23 $T=216660 236640 1 0 $X=216470 $Y=233680
X1213 1 2 ICV_23 $T=216660 258400 1 0 $X=216470 $Y=255440
X1214 1 2 ICV_23 $T=231380 247520 1 0 $X=231190 $Y=244560
X1215 1 2 ICV_23 $T=256220 236640 1 0 $X=256030 $Y=233680
X1216 1 2 ICV_23 $T=272320 242080 0 0 $X=272130 $Y=241840
X1217 1 2 ICV_23 $T=272780 247520 1 0 $X=272590 $Y=244560
X1218 1 2 ICV_23 $T=283820 247520 1 0 $X=283630 $Y=244560
X1219 1 2 ICV_23 $T=286580 247520 0 0 $X=286390 $Y=247280
X1220 1 2 ICV_23 $T=314640 231200 0 0 $X=314450 $Y=230960
X1221 1 2 ICV_23 $T=317400 231200 1 0 $X=317210 $Y=228240
X1222 1 2 ICV_23 $T=319700 225760 0 0 $X=319510 $Y=225520
X1223 1 2 ICV_23 $T=333960 252960 1 0 $X=333770 $Y=250000
X1224 1 2 ICV_24 $T=46460 242080 1 0 $X=46270 $Y=239120
X1225 1 2 ICV_24 $T=46460 263840 1 0 $X=46270 $Y=260880
X1226 1 2 ICV_24 $T=60260 252960 0 0 $X=60070 $Y=252720
X1227 1 2 ICV_24 $T=74520 258400 1 0 $X=74330 $Y=255440
X1228 1 2 ICV_24 $T=102580 225760 1 0 $X=102390 $Y=222800
X1229 1 2 ICV_24 $T=102580 258400 1 0 $X=102390 $Y=255440
X1230 1 2 ICV_24 $T=158700 225760 1 0 $X=158510 $Y=222800
X1231 1 2 ICV_24 $T=172500 247520 0 0 $X=172310 $Y=247280
X1232 1 2 ICV_24 $T=172500 252960 0 0 $X=172310 $Y=252720
X1233 1 2 ICV_24 $T=214820 247520 1 0 $X=214630 $Y=244560
X1234 1 2 ICV_24 $T=214820 263840 1 0 $X=214630 $Y=260880
X1235 1 2 ICV_24 $T=228620 225760 0 0 $X=228430 $Y=225520
X1236 1 2 ICV_24 $T=242880 220320 1 0 $X=242690 $Y=217360
X1237 1 2 ICV_24 $T=270940 225760 1 0 $X=270750 $Y=222800
X1238 1 2 ICV_24 $T=299000 225760 1 0 $X=298810 $Y=222800
X1239 1 2 ICV_24 $T=299000 252960 1 0 $X=298810 $Y=250000
X1240 1 2 ICV_26 $T=5520 220320 0 0 $X=5330 $Y=220080
X1241 1 2 ICV_26 $T=5520 225760 0 0 $X=5330 $Y=225520
X1242 1 2 ICV_26 $T=5520 231200 0 0 $X=5330 $Y=230960
X1243 1 2 ICV_26 $T=5520 236640 0 0 $X=5330 $Y=236400
X1244 1 2 ICV_26 $T=5520 242080 0 0 $X=5330 $Y=241840
X1245 1 2 ICV_26 $T=5520 247520 0 0 $X=5330 $Y=247280
X1246 1 2 ICV_26 $T=5520 252960 0 0 $X=5330 $Y=252720
X1247 1 2 ICV_26 $T=5520 258400 0 0 $X=5330 $Y=258160
X1248 1 2 ICV_26 $T=350520 220320 1 180 $X=348950 $Y=220080
X1249 1 2 ICV_26 $T=350520 225760 1 180 $X=348950 $Y=225520
X1250 1 2 ICV_26 $T=350520 231200 1 180 $X=348950 $Y=230960
X1251 1 2 ICV_26 $T=350520 236640 1 180 $X=348950 $Y=236400
X1252 1 2 ICV_26 $T=350520 242080 1 180 $X=348950 $Y=241840
X1253 1 2 ICV_26 $T=350520 247520 1 180 $X=348950 $Y=247280
X1254 1 2 ICV_26 $T=350520 252960 1 180 $X=348950 $Y=252720
X1255 1 2 ICV_26 $T=350520 258400 1 180 $X=348950 $Y=258160
X1256 1 2 4 376 ICV_27 $T=63020 236640 0 0 $X=62830 $Y=236400
X1257 1 2 43 23 ICV_27 $T=66700 220320 0 0 $X=66510 $Y=220080
X1258 1 2 61 66 ICV_27 $T=71300 220320 1 0 $X=71110 $Y=217360
X1259 1 2 86 87 ICV_27 $T=109480 258400 0 0 $X=109290 $Y=258160
X1260 1 2 4 417 ICV_27 $T=135240 258400 0 0 $X=135050 $Y=258160
X1261 1 2 425 428 ICV_27 $T=161000 231200 0 0 $X=160810 $Y=230960
X1262 1 2 435 441 ICV_27 $T=161460 231200 1 0 $X=161270 $Y=228240
X1263 1 2 442 435 ICV_27 $T=169280 236640 0 0 $X=169090 $Y=236400
X1264 1 2 136 454 ICV_27 $T=180320 242080 0 0 $X=180130 $Y=241840
X1265 1 2 449 456 ICV_27 $T=183080 236640 1 0 $X=182890 $Y=233680
X1266 1 2 466 469 ICV_27 $T=211140 242080 1 0 $X=210950 $Y=239120
X1267 1 2 485 486 ICV_27 $T=239200 252960 1 0 $X=239010 $Y=250000
X1268 1 2 194 498 ICV_27 $T=253460 236640 0 0 $X=253270 $Y=236400
X1269 1 2 499 500 ICV_27 $T=253460 247520 0 0 $X=253270 $Y=247280
X1270 1 2 196 481 ICV_27 $T=253460 258400 0 0 $X=253270 $Y=258160
X1271 1 2 484 486 ICV_27 $T=260360 247520 0 0 $X=260170 $Y=247280
X1272 1 2 530 196 ICV_27 $T=309580 242080 0 0 $X=309390 $Y=241840
X1273 1 2 236 350 ICV_27 $T=316020 225760 1 0 $X=315830 $Y=222800
X1274 1 2 3 4 ICV_27 $T=337180 258400 0 0 $X=336990 $Y=258160
X1275 1 2 43 ICV_28 $T=58880 220320 0 0 $X=58690 $Y=220080
X1276 1 2 64 ICV_28 $T=73140 225760 1 0 $X=72950 $Y=222800
X1277 1 2 49 ICV_28 $T=86940 225760 0 0 $X=86750 $Y=225520
X1278 1 2 393 ICV_28 $T=101200 252960 1 0 $X=101010 $Y=250000
X1279 1 2 89 ICV_28 $T=115000 225760 0 0 $X=114810 $Y=225520
X1280 1 2 114 ICV_28 $T=143060 231200 0 0 $X=142870 $Y=230960
X1281 1 2 419 ICV_28 $T=143060 242080 0 0 $X=142870 $Y=241840
X1282 1 2 131 ICV_28 $T=171120 242080 0 0 $X=170930 $Y=241840
X1283 1 2 455 ICV_28 $T=199180 225760 0 0 $X=198990 $Y=225520
X1284 1 2 178 ICV_28 $T=227240 220320 0 0 $X=227050 $Y=220080
X1285 1 2 136 ICV_28 $T=227240 247520 0 0 $X=227050 $Y=247280
X1286 1 2 487 ICV_28 $T=241500 258400 1 0 $X=241310 $Y=255440
X1287 1 2 486 ICV_28 $T=255300 242080 0 0 $X=255110 $Y=241840
X1288 1 2 172 ICV_28 $T=283360 231200 0 0 $X=283170 $Y=230960
X1289 1 2 227 ICV_28 $T=311420 220320 0 0 $X=311230 $Y=220080
X1290 1 2 524 ICV_28 $T=311420 225760 0 0 $X=311230 $Y=225520
X1291 1 2 235 ICV_28 $T=311420 231200 0 0 $X=311230 $Y=230960
X1292 1 2 526 ICV_28 $T=311420 247520 0 0 $X=311230 $Y=247280
X1293 1 2 526 ICV_28 $T=311420 252960 0 0 $X=311230 $Y=252720
X1294 1 2 535 ICV_28 $T=325680 258400 1 0 $X=325490 $Y=255440
X1295 1 2 ICV_29 $T=10580 220320 1 0 $X=10390 $Y=217360
X1296 1 2 ICV_29 $T=10580 231200 1 0 $X=10390 $Y=228240
X1297 1 2 ICV_29 $T=10580 242080 1 0 $X=10390 $Y=239120
X1298 1 2 ICV_29 $T=10580 247520 1 0 $X=10390 $Y=244560
X1299 1 2 ICV_29 $T=10580 252960 1 0 $X=10390 $Y=250000
X1300 1 2 ICV_29 $T=23920 258400 0 0 $X=23730 $Y=258160
X1301 1 2 ICV_29 $T=38640 252960 1 0 $X=38450 $Y=250000
X1302 1 2 ICV_29 $T=46460 252960 0 0 $X=46270 $Y=252720
X1303 1 2 ICV_29 $T=57040 258400 1 0 $X=56850 $Y=255440
X1304 1 2 ICV_29 $T=83720 236640 1 0 $X=83530 $Y=233680
X1305 1 2 ICV_29 $T=88320 247520 1 0 $X=88130 $Y=244560
X1306 1 2 ICV_29 $T=104420 225760 1 0 $X=104230 $Y=222800
X1307 1 2 ICV_29 $T=133860 225760 0 0 $X=133670 $Y=225520
X1308 1 2 ICV_29 $T=135700 247520 0 0 $X=135510 $Y=247280
X1309 1 2 ICV_29 $T=137540 220320 1 0 $X=137350 $Y=217360
X1310 1 2 ICV_29 $T=162840 220320 0 0 $X=162650 $Y=220080
X1311 1 2 ICV_29 $T=164680 225760 0 0 $X=164490 $Y=225520
X1312 1 2 ICV_29 $T=195040 263840 1 0 $X=194850 $Y=260880
X1313 1 2 ICV_29 $T=195960 242080 1 0 $X=195770 $Y=239120
X1314 1 2 ICV_29 $T=216660 231200 1 0 $X=216470 $Y=228240
X1315 1 2 ICV_29 $T=230460 247520 0 0 $X=230270 $Y=247280
X1316 1 2 ICV_29 $T=258520 236640 0 0 $X=258330 $Y=236400
X1317 1 2 ICV_29 $T=262660 242080 1 0 $X=262470 $Y=239120
X1318 1 2 ICV_29 $T=263120 231200 1 0 $X=262930 $Y=228240
X1319 1 2 ICV_29 $T=290260 258400 0 0 $X=290070 $Y=258160
X1320 1 2 ICV_29 $T=290720 263840 1 0 $X=290530 $Y=260880
X1321 1 2 ICV_29 $T=318780 263840 1 0 $X=318590 $Y=260880
X1322 1 2 13 13 17 354 ICV_30 $T=21160 220320 0 0 $X=20970 $Y=220080
X1323 1 2 361 15 361 359 ICV_30 $T=26220 242080 1 0 $X=26030 $Y=239120
X1324 1 2 40 40 41 375 ICV_30 $T=51060 258400 0 0 $X=50870 $Y=258160
X1325 1 2 58 58 380 378 ICV_30 $T=67620 242080 0 0 $X=67430 $Y=241840
X1326 1 2 15 15 383 67 ICV_30 $T=69000 225760 0 0 $X=68810 $Y=225520
X1327 1 2 75 75 397 394 ICV_30 $T=93380 242080 0 0 $X=93190 $Y=241840
X1328 1 2 85 86 87 406 ICV_30 $T=105340 263840 1 0 $X=105150 $Y=260880
X1329 1 2 403 88 403 399 ICV_30 $T=108100 220320 0 0 $X=107910 $Y=220080
X1330 1 2 409 75 408 413 ICV_30 $T=118220 252960 1 0 $X=118030 $Y=250000
X1331 1 2 418 109 419 415 ICV_30 $T=136620 247520 1 0 $X=136430 $Y=244560
X1332 1 2 430 109 430 436 ICV_30 $T=150420 258400 1 0 $X=150230 $Y=255440
X1333 1 2 162 161 463 165 ICV_30 $T=205160 263840 1 0 $X=204970 $Y=260880
X1334 1 2 161 161 471 476 ICV_30 $T=217120 242080 0 0 $X=216930 $Y=241840
X1335 1 2 164 164 475 477 ICV_30 $T=220340 220320 0 0 $X=220150 $Y=220080
X1336 1 2 185 185 490 491 ICV_30 $T=242880 220320 0 0 $X=242690 $Y=220080
X1337 1 2 189 184 493 489 ICV_30 $T=245640 247520 1 0 $X=245450 $Y=244560
X1338 1 2 481 184 502 505 ICV_30 $T=262660 258400 1 0 $X=262470 $Y=255440
X1339 1 2 184 184 503 506 ICV_30 $T=262660 258400 0 0 $X=262470 $Y=258160
.ENDS
***************************************
.SUBCKT ICV_32 1 2
** N=2 EP=2 IP=4 FDC=4
*.SEEDPROM
X1 1 2 ICV_23 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269
** N=586 EP=269 IP=5674 FDC=7968
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=178105 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=183545 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=188985 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=194425 $D=191
X4 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=199865 $D=191
X5 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=205305 $D=191
X6 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=210745 $D=191
X7 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=8740 182240 1 0 $X=8550 $Y=179280
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=22080 193120 1 0 $X=21890 $Y=190160
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=32660 176800 1 0 $X=32470 $Y=173840
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=46460 193120 1 0 $X=46270 $Y=190160
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=46460 214880 1 0 $X=46270 $Y=211920
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=48760 193120 0 0 $X=48570 $Y=192880
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=53820 209440 1 0 $X=53630 $Y=206480
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=55200 198560 0 0 $X=55010 $Y=198320
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=58420 176800 0 0 $X=58230 $Y=176560
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=58420 214880 0 0 $X=58230 $Y=214640
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=62100 193120 0 0 $X=61910 $Y=192880
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74520 209440 1 0 $X=74330 $Y=206480
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 214880 0 0 $X=76170 $Y=214640
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=80500 214880 0 0 $X=80310 $Y=214640
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=84640 204000 0 0 $X=84450 $Y=203760
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=86480 209440 0 0 $X=86290 $Y=209200
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88320 214880 0 0 $X=88130 $Y=214640
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=91080 209440 1 0 $X=90890 $Y=206480
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=97520 182240 1 0 $X=97330 $Y=179280
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 187680 1 0 $X=102390 $Y=184720
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=116380 209440 0 0 $X=116190 $Y=209200
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 198560 0 0 $X=118030 $Y=198320
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 209440 0 0 $X=118030 $Y=209200
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118680 214880 1 0 $X=118490 $Y=211920
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=120520 209440 1 0 $X=120330 $Y=206480
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=122820 182240 1 0 $X=122630 $Y=179280
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=127880 176800 0 0 $X=127690 $Y=176560
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 204000 1 0 $X=130450 $Y=201040
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=142600 182240 0 0 $X=142410 $Y=182000
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 193120 0 0 $X=144250 $Y=192880
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=146280 176800 0 0 $X=146090 $Y=176560
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 187680 1 0 $X=158510 $Y=184720
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 193120 1 0 $X=158510 $Y=190160
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 176800 1 0 $X=160350 $Y=173840
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 214880 1 0 $X=160350 $Y=211920
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 214880 0 0 $X=174150 $Y=214640
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=178940 176800 1 0 $X=178750 $Y=173840
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=192280 209440 0 0 $X=192090 $Y=209200
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=192280 214880 1 0 $X=192090 $Y=211920
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=195960 182240 1 0 $X=195770 $Y=179280
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=199640 204000 1 0 $X=199450 $Y=201040
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 182240 1 0 $X=202210 $Y=179280
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=203320 193120 1 0 $X=203130 $Y=190160
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=209300 214880 0 0 $X=209110 $Y=214640
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=212980 209440 1 0 $X=212790 $Y=206480
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 198560 1 0 $X=214630 $Y=195600
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220340 198560 1 0 $X=220150 $Y=195600
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=223100 193120 0 0 $X=222910 $Y=192880
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224940 176800 0 0 $X=224750 $Y=176560
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=232300 176800 0 0 $X=232110 $Y=176560
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=235980 176800 1 0 $X=235790 $Y=173840
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 187680 1 0 $X=242690 $Y=184720
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=243800 214880 0 0 $X=243610 $Y=214640
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=244260 182240 0 0 $X=244070 $Y=182000
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=253460 209440 0 0 $X=253270 $Y=209200
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=256680 182240 0 0 $X=256490 $Y=182000
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=264040 187680 0 0 $X=263850 $Y=187440
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 176800 1 0 $X=270750 $Y=173840
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=275540 193120 0 0 $X=275350 $Y=192880
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 182240 0 0 $X=284550 $Y=182000
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286580 198560 0 0 $X=286390 $Y=198320
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=287500 176800 1 0 $X=287310 $Y=173840
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=288420 214880 0 0 $X=288230 $Y=214640
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=297160 193120 1 0 $X=296970 $Y=190160
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 182240 1 0 $X=298810 $Y=179280
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 198560 1 0 $X=298810 $Y=195600
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 204000 1 0 $X=298810 $Y=201040
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 209440 1 0 $X=300650 $Y=206480
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=306360 204000 1 0 $X=306170 $Y=201040
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=309120 176800 0 0 $X=308930 $Y=176560
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=309120 209440 1 0 $X=308930 $Y=206480
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=309120 214880 1 0 $X=308930 $Y=211920
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=327060 193120 1 0 $X=326870 $Y=190160
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=332580 176800 1 0 $X=332390 $Y=173840
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=332580 182240 1 0 $X=332390 $Y=179280
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=332580 187680 1 0 $X=332390 $Y=184720
X83 1 2 ICV_1 $T=5520 176800 1 0 $X=5330 $Y=173840
X84 1 2 ICV_1 $T=5520 182240 1 0 $X=5330 $Y=179280
X85 1 2 ICV_1 $T=5520 187680 1 0 $X=5330 $Y=184720
X86 1 2 ICV_1 $T=5520 193120 1 0 $X=5330 $Y=190160
X87 1 2 ICV_1 $T=5520 198560 1 0 $X=5330 $Y=195600
X88 1 2 ICV_1 $T=5520 204000 1 0 $X=5330 $Y=201040
X89 1 2 ICV_1 $T=5520 209440 1 0 $X=5330 $Y=206480
X90 1 2 ICV_1 $T=5520 214880 1 0 $X=5330 $Y=211920
X91 1 2 ICV_1 $T=350520 176800 0 180 $X=348950 $Y=173840
X92 1 2 ICV_1 $T=350520 182240 0 180 $X=348950 $Y=179280
X93 1 2 ICV_1 $T=350520 187680 0 180 $X=348950 $Y=184720
X94 1 2 ICV_1 $T=350520 193120 0 180 $X=348950 $Y=190160
X95 1 2 ICV_1 $T=350520 198560 0 180 $X=348950 $Y=195600
X96 1 2 ICV_1 $T=350520 204000 0 180 $X=348950 $Y=201040
X97 1 2 ICV_1 $T=350520 209440 0 180 $X=348950 $Y=206480
X98 1 2 ICV_1 $T=350520 214880 0 180 $X=348950 $Y=211920
X194 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=24380 187680 1 0 $X=24190 $Y=184720
X195 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=28980 176800 1 0 $X=28790 $Y=173840
X196 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 176800 1 0 $X=43970 $Y=173840
X197 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 182240 1 0 $X=43970 $Y=179280
X198 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 209440 1 0 $X=43970 $Y=206480
X199 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=50600 187680 1 0 $X=50410 $Y=184720
X200 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=51520 182240 0 0 $X=51330 $Y=182000
X201 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=54740 214880 0 0 $X=54550 $Y=214640
X202 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 182240 0 0 $X=57770 $Y=182000
X203 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=58420 193120 1 0 $X=58230 $Y=190160
X204 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=60720 198560 1 0 $X=60530 $Y=195600
X205 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=62100 198560 0 0 $X=61910 $Y=198320
X206 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=68540 198560 1 0 $X=68350 $Y=195600
X207 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71760 198560 0 0 $X=71570 $Y=198320
X208 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 176800 1 0 $X=72030 $Y=173840
X209 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 204000 1 0 $X=76170 $Y=201040
X210 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=86940 182240 1 0 $X=86750 $Y=179280
X211 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 182240 1 0 $X=100090 $Y=179280
X212 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=109480 209440 1 0 $X=109290 $Y=206480
X213 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=113620 176800 0 0 $X=113430 $Y=176560
X214 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=136620 182240 0 0 $X=136430 $Y=182000
X215 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=138000 187680 1 0 $X=137810 $Y=184720
X216 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 176800 1 0 $X=139650 $Y=173840
X217 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=143520 204000 1 0 $X=143330 $Y=201040
X218 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=155020 193120 1 0 $X=154830 $Y=190160
X219 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=155480 209440 1 0 $X=155290 $Y=206480
X220 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 204000 1 0 $X=156210 $Y=201040
X221 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=157320 209440 0 0 $X=157130 $Y=209200
X222 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=159160 187680 0 0 $X=158970 $Y=187440
X223 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=159160 193120 0 0 $X=158970 $Y=192880
X224 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=166060 204000 0 0 $X=165870 $Y=203760
X225 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=172500 182240 1 0 $X=172310 $Y=179280
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=179400 204000 0 0 $X=179210 $Y=203760
X227 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184000 204000 1 0 $X=183810 $Y=201040
X228 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 187680 0 0 $X=184270 $Y=187440
X229 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 209440 1 0 $X=184270 $Y=206480
X230 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 214880 1 0 $X=188410 $Y=211920
X231 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=190900 193120 1 0 $X=190710 $Y=190160
X232 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=190900 198560 1 0 $X=190710 $Y=195600
X233 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198260 204000 0 0 $X=198070 $Y=203760
X234 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198720 182240 1 0 $X=198530 $Y=179280
X235 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=201940 176800 1 0 $X=201750 $Y=173840
X236 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=207000 176800 1 0 $X=206810 $Y=173840
X237 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 198560 1 0 $X=210950 $Y=195600
X238 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212060 187680 1 0 $X=211870 $Y=184720
X239 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 198560 1 0 $X=216470 $Y=195600
X240 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=217120 214880 0 0 $X=216930 $Y=214640
X241 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=221720 176800 1 0 $X=221530 $Y=173840
X242 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=223100 214880 1 0 $X=222910 $Y=211920
X243 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 182240 0 0 $X=226130 $Y=182000
X244 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 187680 0 0 $X=230270 $Y=187440
X245 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=232300 176800 1 0 $X=232110 $Y=173840
X246 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=235980 214880 0 0 $X=235790 $Y=214640
X247 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239200 187680 1 0 $X=239010 $Y=184720
X248 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239660 198560 1 0 $X=239470 $Y=195600
X249 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=251160 214880 1 0 $X=250970 $Y=211920
X250 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=253000 182240 0 0 $X=252810 $Y=182000
X251 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254380 204000 1 0 $X=254190 $Y=201040
X252 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254840 198560 1 0 $X=254650 $Y=195600
X253 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=261280 214880 1 0 $X=261090 $Y=211920
X254 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=262660 182240 1 0 $X=262470 $Y=179280
X255 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=263120 209440 1 0 $X=262930 $Y=206480
X256 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=266340 214880 1 0 $X=266150 $Y=211920
X257 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267260 176800 1 0 $X=267070 $Y=173840
X258 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 204000 1 0 $X=268450 $Y=201040
X259 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278300 209440 0 0 $X=278110 $Y=209200
X260 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=280140 209440 1 0 $X=279950 $Y=206480
X261 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281520 198560 0 0 $X=281330 $Y=198320
X262 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=283820 176800 1 0 $X=283630 $Y=173840
X263 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286580 193120 0 0 $X=286390 $Y=192880
X264 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 209440 1 0 $X=296510 $Y=206480
X265 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 214880 1 0 $X=296510 $Y=211920
X266 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=303600 198560 0 0 $X=303410 $Y=198320
X267 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=306360 198560 1 0 $X=306170 $Y=195600
X268 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=308660 204000 0 0 $X=308470 $Y=203760
X269 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 198560 1 0 $X=324570 $Y=195600
X270 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 204000 1 0 $X=324570 $Y=201040
X271 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 176800 1 0 $X=328710 $Y=173840
X272 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 182240 1 0 $X=328710 $Y=179280
X273 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 187680 1 0 $X=328710 $Y=184720
X274 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=337640 209440 0 0 $X=337450 $Y=209200
X275 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344540 176800 1 0 $X=344350 $Y=173840
X276 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344540 182240 1 0 $X=344350 $Y=179280
X277 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344540 187680 1 0 $X=344350 $Y=184720
X278 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 193120 1 0 $X=344810 $Y=190160
X279 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 198560 1 0 $X=345270 $Y=195600
X280 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 204000 1 0 $X=345270 $Y=201040
X281 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=20700 182240 0 0 $X=20510 $Y=182000
X282 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25300 182240 1 0 $X=25110 $Y=179280
X283 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40940 214880 1 0 $X=40750 $Y=211920
X284 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=48300 204000 1 0 $X=48110 $Y=201040
X285 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55660 214880 1 0 $X=55470 $Y=211920
X286 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=60720 209440 1 0 $X=60530 $Y=206480
X287 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=63480 182240 1 0 $X=63290 $Y=179280
X288 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=67160 204000 1 0 $X=66970 $Y=201040
X289 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=70840 187680 0 0 $X=70650 $Y=187440
X290 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=73140 182240 0 0 $X=72950 $Y=182000
X291 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=79120 204000 0 0 $X=78930 $Y=203760
X292 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81880 204000 1 0 $X=81690 $Y=201040
X293 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82800 193120 1 0 $X=82610 $Y=190160
X294 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=92000 182240 1 0 $X=91810 $Y=179280
X295 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=96600 176800 1 0 $X=96410 $Y=173840
X296 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=110860 198560 1 0 $X=110670 $Y=195600
X297 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=112240 187680 0 0 $X=112050 $Y=187440
X298 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 182240 1 0 $X=125390 $Y=179280
X299 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=126500 187680 1 0 $X=126310 $Y=184720
X300 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=137540 187680 0 0 $X=137350 $Y=187440
X301 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=138920 193120 0 0 $X=138730 $Y=192880
X302 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=159620 176800 0 0 $X=159430 $Y=176560
X303 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=163300 198560 0 0 $X=163110 $Y=198320
X304 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=182620 198560 1 0 $X=182430 $Y=195600
X305 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=196420 193120 1 0 $X=196230 $Y=190160
X306 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=196420 198560 1 0 $X=196230 $Y=195600
X307 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=196420 209440 0 0 $X=196230 $Y=209200
X308 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=199640 187680 1 0 $X=199450 $Y=184720
X309 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=202400 204000 1 0 $X=202210 $Y=201040
X310 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=208840 193120 1 0 $X=208650 $Y=190160
X311 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210220 182240 1 0 $X=210030 $Y=179280
X312 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=222180 187680 0 0 $X=221990 $Y=187440
X313 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=231840 182240 1 0 $X=231650 $Y=179280
X314 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=236440 214880 1 0 $X=236250 $Y=211920
X315 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=238740 193120 1 0 $X=238550 $Y=190160
X316 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=241960 193120 0 0 $X=241770 $Y=192880
X317 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=250700 198560 0 0 $X=250510 $Y=198320
X318 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=262200 214880 0 0 $X=262010 $Y=214640
X319 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=280140 204000 0 0 $X=279950 $Y=203760
X320 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=295320 214880 0 0 $X=295130 $Y=214640
X321 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=305900 187680 1 0 $X=305710 $Y=184720
X322 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=307280 182240 1 0 $X=307090 $Y=179280
X323 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=308200 182240 0 0 $X=308010 $Y=182000
X324 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=319240 193120 1 0 $X=319050 $Y=190160
X325 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=325680 182240 0 0 $X=325490 $Y=182000
X326 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=326140 176800 0 0 $X=325950 $Y=176560
X327 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=326140 187680 0 0 $X=325950 $Y=187440
X328 1 2 ICV_2 $T=75900 182240 1 0 $X=75710 $Y=179280
X329 1 2 ICV_2 $T=132020 187680 1 0 $X=131830 $Y=184720
X330 1 2 ICV_2 $T=145820 198560 0 0 $X=145630 $Y=198320
X331 1 2 ICV_2 $T=160080 193120 1 0 $X=159890 $Y=190160
X332 1 2 ICV_2 $T=160080 198560 1 0 $X=159890 $Y=195600
X333 1 2 ICV_2 $T=201940 176800 0 0 $X=201750 $Y=176560
X334 1 2 ICV_2 $T=230000 182240 0 0 $X=229810 $Y=182000
X335 1 2 ICV_2 $T=230000 214880 0 0 $X=229810 $Y=214640
X336 1 2 ICV_2 $T=258060 182240 0 0 $X=257870 $Y=182000
X337 1 2 ICV_2 $T=258060 187680 0 0 $X=257870 $Y=187440
X338 1 2 ICV_2 $T=300380 176800 1 0 $X=300190 $Y=173840
X339 1 2 ICV_2 $T=300380 198560 1 0 $X=300190 $Y=195600
X340 1 2 ICV_2 $T=300380 204000 1 0 $X=300190 $Y=201040
X341 1 2 ICV_2 $T=328440 193120 1 0 $X=328250 $Y=190160
X342 1 2 ICV_2 $T=328440 198560 1 0 $X=328250 $Y=195600
X343 1 2 ICV_2 $T=328440 204000 1 0 $X=328250 $Y=201040
X344 1 2 ICV_2 $T=328440 214880 1 0 $X=328250 $Y=211920
X345 1 2 ICV_2 $T=342240 176800 0 0 $X=342050 $Y=176560
X346 1 2 ICV_2 $T=342240 182240 0 0 $X=342050 $Y=182000
X347 1 2 ICV_2 $T=342240 187680 0 0 $X=342050 $Y=187440
X348 1 2 ICV_2 $T=342240 198560 0 0 $X=342050 $Y=198320
X349 1 2 ICV_2 $T=342240 204000 0 0 $X=342050 $Y=203760
X350 1 2 ICV_2 $T=342240 209440 0 0 $X=342050 $Y=209200
X351 1 2 ICV_2 $T=342240 214880 0 0 $X=342050 $Y=214640
X352 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 187680 1 0 $X=17750 $Y=184720
X353 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 193120 1 0 $X=17750 $Y=190160
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 193120 0 0 $X=18210 $Y=192880
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 209440 0 0 $X=18210 $Y=209200
X356 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=25300 187680 0 0 $X=25110 $Y=187440
X357 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=27600 214880 0 0 $X=27410 $Y=214640
X358 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 198560 1 0 $X=31550 $Y=195600
X359 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=48300 198560 1 0 $X=48110 $Y=195600
X360 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=51980 193120 1 0 $X=51790 $Y=190160
X361 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=61180 214880 1 0 $X=60990 $Y=211920
X362 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=65780 176800 1 0 $X=65590 $Y=173840
X363 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69000 182240 1 0 $X=68810 $Y=179280
X364 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=85560 198560 1 0 $X=85370 $Y=195600
X365 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=96600 204000 1 0 $X=96410 $Y=201040
X366 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=96600 209440 1 0 $X=96410 $Y=206480
X367 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=101660 214880 1 0 $X=101470 $Y=211920
X368 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 176800 1 0 $X=101930 $Y=173840
X369 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=109020 198560 0 0 $X=108830 $Y=198320
X370 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=111780 204000 0 0 $X=111590 $Y=203760
X371 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 182240 1 0 $X=115730 $Y=179280
X372 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=121440 176800 1 0 $X=121250 $Y=173840
X373 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=130180 193120 1 0 $X=129990 $Y=190160
X374 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 198560 1 0 $X=143330 $Y=195600
X375 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=153180 176800 1 0 $X=152990 $Y=173840
X376 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=157780 198560 1 0 $X=157590 $Y=195600
X377 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158700 198560 0 0 $X=158510 $Y=198320
X378 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172500 176800 1 0 $X=172310 $Y=173840
X379 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=189520 204000 0 0 $X=189330 $Y=203760
X380 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=203320 198560 1 0 $X=203130 $Y=195600
X381 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 193120 1 0 $X=214170 $Y=190160
X382 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=227700 187680 0 0 $X=227510 $Y=187440
X383 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=228160 214880 1 0 $X=227970 $Y=211920
X384 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=235980 182240 0 0 $X=235790 $Y=182000
X385 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244720 209440 1 0 $X=244530 $Y=206480
X386 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=256220 198560 0 0 $X=256030 $Y=198320
X387 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=272780 193120 1 0 $X=272590 $Y=190160
X388 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286580 182240 1 0 $X=286390 $Y=179280
X389 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286580 193120 1 0 $X=286390 $Y=190160
X390 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=303140 214880 1 0 $X=302950 $Y=211920
X391 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=308660 193120 0 0 $X=308470 $Y=192880
X392 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=331660 176800 0 0 $X=331470 $Y=176560
X393 1 4 sky130_fd_sc_hd__diode_2 $T=7820 182240 1 0 $X=7630 $Y=179280
X394 1 4 sky130_fd_sc_hd__diode_2 $T=7820 204000 1 0 $X=7630 $Y=201040
X395 1 370 sky130_fd_sc_hd__diode_2 $T=7820 204000 0 0 $X=7630 $Y=203760
X396 1 13 sky130_fd_sc_hd__diode_2 $T=19320 176800 0 0 $X=19130 $Y=176560
X397 1 14 sky130_fd_sc_hd__diode_2 $T=19320 187680 0 0 $X=19130 $Y=187440
X398 1 373 sky130_fd_sc_hd__diode_2 $T=19320 198560 0 0 $X=19130 $Y=198320
X399 1 375 sky130_fd_sc_hd__diode_2 $T=21160 187680 1 0 $X=20970 $Y=184720
X400 1 376 sky130_fd_sc_hd__diode_2 $T=21160 193120 1 0 $X=20970 $Y=190160
X401 1 370 sky130_fd_sc_hd__diode_2 $T=21620 214880 0 0 $X=21430 $Y=214640
X402 1 382 sky130_fd_sc_hd__diode_2 $T=31740 209440 1 0 $X=31550 $Y=206480
X403 1 27 sky130_fd_sc_hd__diode_2 $T=32660 214880 1 0 $X=32470 $Y=211920
X404 1 28 sky130_fd_sc_hd__diode_2 $T=34040 198560 1 0 $X=33850 $Y=195600
X405 1 36 sky130_fd_sc_hd__diode_2 $T=40020 204000 0 0 $X=39830 $Y=203760
X406 1 37 sky130_fd_sc_hd__diode_2 $T=41400 193120 0 0 $X=41210 $Y=192880
X407 1 396 sky130_fd_sc_hd__diode_2 $T=45080 214880 0 0 $X=44890 $Y=214640
X408 1 40 sky130_fd_sc_hd__diode_2 $T=47840 187680 0 0 $X=47650 $Y=187440
X409 1 401 sky130_fd_sc_hd__diode_2 $T=54280 198560 0 0 $X=54090 $Y=198320
X410 1 58 sky130_fd_sc_hd__diode_2 $T=65780 198560 0 0 $X=65590 $Y=198320
X411 1 4 sky130_fd_sc_hd__diode_2 $T=69460 176800 0 0 $X=69270 $Y=176560
X412 1 66 sky130_fd_sc_hd__diode_2 $T=75440 214880 0 0 $X=75250 $Y=214640
X413 1 68 sky130_fd_sc_hd__diode_2 $T=77280 176800 1 0 $X=77090 $Y=173840
X414 1 52 sky130_fd_sc_hd__diode_2 $T=78200 198560 0 0 $X=78010 $Y=198320
X415 1 76 sky130_fd_sc_hd__diode_2 $T=85560 209440 0 0 $X=85370 $Y=209200
X416 1 416 sky130_fd_sc_hd__diode_2 $T=88320 193120 1 0 $X=88130 $Y=190160
X417 1 417 sky130_fd_sc_hd__diode_2 $T=88320 204000 1 0 $X=88130 $Y=201040
X418 1 418 sky130_fd_sc_hd__diode_2 $T=90160 209440 1 0 $X=89970 $Y=206480
X419 1 4 sky130_fd_sc_hd__diode_2 $T=93380 214880 0 0 $X=93190 $Y=214640
X420 1 422 sky130_fd_sc_hd__diode_2 $T=94760 193120 0 0 $X=94570 $Y=192880
X421 1 83 sky130_fd_sc_hd__diode_2 $T=97060 204000 0 0 $X=96870 $Y=203760
X422 1 80 sky130_fd_sc_hd__diode_2 $T=100280 187680 0 0 $X=100090 $Y=187440
X423 1 52 sky130_fd_sc_hd__diode_2 $T=100740 182240 0 0 $X=100550 $Y=182000
X424 1 404 sky130_fd_sc_hd__diode_2 $T=109020 193120 1 0 $X=108830 $Y=190160
X425 1 89 sky130_fd_sc_hd__diode_2 $T=109480 176800 1 0 $X=109290 $Y=173840
X426 1 103 sky130_fd_sc_hd__diode_2 $T=130640 182240 0 0 $X=130450 $Y=182000
X427 1 95 sky130_fd_sc_hd__diode_2 $T=132020 214880 0 0 $X=131830 $Y=214640
X428 1 439 sky130_fd_sc_hd__diode_2 $T=134780 209440 0 0 $X=134590 $Y=209200
X429 1 442 sky130_fd_sc_hd__diode_2 $T=143980 182240 1 0 $X=143790 $Y=179280
X430 1 443 sky130_fd_sc_hd__diode_2 $T=144900 214880 1 0 $X=144710 $Y=211920
X431 1 120 sky130_fd_sc_hd__diode_2 $T=147200 193120 0 0 $X=147010 $Y=192880
X432 1 4 sky130_fd_sc_hd__diode_2 $T=148120 204000 1 0 $X=147930 $Y=201040
X433 1 122 sky130_fd_sc_hd__diode_2 $T=152260 214880 0 0 $X=152070 $Y=214640
X434 1 4 sky130_fd_sc_hd__diode_2 $T=158700 182240 0 0 $X=158510 $Y=182000
X435 1 459 sky130_fd_sc_hd__diode_2 $T=172960 187680 1 0 $X=172770 $Y=184720
X436 1 139 sky130_fd_sc_hd__diode_2 $T=173420 193120 1 0 $X=173230 $Y=190160
X437 1 464 sky130_fd_sc_hd__diode_2 $T=174340 198560 1 0 $X=174150 $Y=195600
X438 1 4 sky130_fd_sc_hd__diode_2 $T=175720 214880 1 0 $X=175530 $Y=211920
X439 1 465 sky130_fd_sc_hd__diode_2 $T=176180 182240 1 0 $X=175990 $Y=179280
X440 1 460 sky130_fd_sc_hd__diode_2 $T=178020 176800 1 0 $X=177830 $Y=173840
X441 1 143 sky130_fd_sc_hd__diode_2 $T=180320 182240 0 0 $X=180130 $Y=182000
X442 1 151 sky130_fd_sc_hd__diode_2 $T=188140 187680 0 0 $X=187950 $Y=187440
X443 1 468 sky130_fd_sc_hd__diode_2 $T=202400 193120 1 0 $X=202210 $Y=190160
X444 1 4 sky130_fd_sc_hd__diode_2 $T=203320 198560 0 0 $X=203130 $Y=198320
X445 1 175 sky130_fd_sc_hd__diode_2 $T=204700 182240 0 0 $X=204510 $Y=182000
X446 1 97 sky130_fd_sc_hd__diode_2 $T=208380 214880 0 0 $X=208190 $Y=214640
X447 1 4 sky130_fd_sc_hd__diode_2 $T=208840 176800 0 0 $X=208650 $Y=176560
X448 1 179 sky130_fd_sc_hd__diode_2 $T=210680 204000 0 0 $X=210490 $Y=203760
X449 1 178 sky130_fd_sc_hd__diode_2 $T=220340 198560 0 0 $X=220150 $Y=198320
X450 1 186 sky130_fd_sc_hd__diode_2 $T=224940 209440 1 0 $X=224750 $Y=206480
X451 1 116 sky130_fd_sc_hd__diode_2 $T=231380 176800 0 0 $X=231190 $Y=176560
X452 1 198 sky130_fd_sc_hd__diode_2 $T=234600 187680 0 0 $X=234410 $Y=187440
X453 1 487 sky130_fd_sc_hd__diode_2 $T=238280 182240 0 0 $X=238090 $Y=182000
X454 1 122 sky130_fd_sc_hd__diode_2 $T=242880 214880 0 0 $X=242690 $Y=214640
X455 1 186 sky130_fd_sc_hd__diode_2 $T=245180 209440 0 0 $X=244990 $Y=209200
X456 1 203 sky130_fd_sc_hd__diode_2 $T=247020 209440 1 0 $X=246830 $Y=206480
X457 1 217 sky130_fd_sc_hd__diode_2 $T=263120 204000 0 0 $X=262930 $Y=203760
X458 1 4 sky130_fd_sc_hd__diode_2 $T=264960 182240 0 0 $X=264770 $Y=182000
X459 1 219 sky130_fd_sc_hd__diode_2 $T=268640 214880 0 0 $X=268450 $Y=214640
X460 1 222 sky130_fd_sc_hd__diode_2 $T=272780 214880 0 0 $X=272590 $Y=214640
X461 1 504 sky130_fd_sc_hd__diode_2 $T=274620 193120 0 0 $X=274430 $Y=192880
X462 1 508 sky130_fd_sc_hd__diode_2 $T=286120 187680 1 0 $X=285930 $Y=184720
X463 1 230 sky130_fd_sc_hd__diode_2 $T=287500 182240 0 0 $X=287310 $Y=182000
X464 1 226 sky130_fd_sc_hd__diode_2 $T=287500 214880 0 0 $X=287310 $Y=214640
X465 1 4 sky130_fd_sc_hd__diode_2 $T=288880 204000 0 0 $X=288690 $Y=203760
X466 1 516 sky130_fd_sc_hd__diode_2 $T=290720 209440 1 0 $X=290530 $Y=206480
X467 1 517 sky130_fd_sc_hd__diode_2 $T=291640 198560 0 0 $X=291450 $Y=198320
X468 1 515 sky130_fd_sc_hd__diode_2 $T=292100 182240 1 0 $X=291910 $Y=179280
X469 1 251 sky130_fd_sc_hd__diode_2 $T=306360 176800 1 0 $X=306170 $Y=173840
X470 1 253 sky130_fd_sc_hd__diode_2 $T=308200 214880 1 0 $X=308010 $Y=211920
X471 1 257 sky130_fd_sc_hd__diode_2 $T=312800 182240 1 0 $X=312610 $Y=179280
X472 1 4 sky130_fd_sc_hd__diode_2 $T=324300 193120 0 0 $X=324110 $Y=192880
X473 1 534 sky130_fd_sc_hd__diode_2 $T=325680 209440 0 0 $X=325490 $Y=209200
X474 1 2 4 ICV_4 $T=20240 193120 0 0 $X=20050 $Y=192880
X475 1 2 4 ICV_4 $T=20240 209440 0 0 $X=20050 $Y=209200
X476 1 2 20 ICV_4 $T=35880 187680 1 0 $X=35690 $Y=184720
X477 1 2 390 ICV_4 $T=38640 193120 1 0 $X=38450 $Y=190160
X478 1 2 34 ICV_4 $T=40020 176800 0 0 $X=39830 $Y=176560
X479 1 2 390 ICV_4 $T=42320 214880 0 0 $X=42130 $Y=214640
X480 1 2 33 ICV_4 $T=43240 182240 0 0 $X=43050 $Y=182000
X481 1 2 24 ICV_4 $T=43240 198560 1 0 $X=43050 $Y=195600
X482 1 2 43 ICV_4 $T=51980 187680 0 0 $X=51790 $Y=187440
X483 1 2 23 ICV_4 $T=54280 193120 1 0 $X=54090 $Y=190160
X484 1 2 404 ICV_4 $T=58880 204000 0 0 $X=58690 $Y=203760
X485 1 2 39 ICV_4 $T=58880 209440 0 0 $X=58690 $Y=209200
X486 1 2 26 ICV_4 $T=65320 214880 0 0 $X=65130 $Y=214640
X487 1 2 400 ICV_4 $T=69920 193120 0 0 $X=69730 $Y=192880
X488 1 2 64 ICV_4 $T=73140 193120 1 0 $X=72950 $Y=190160
X489 1 2 65 ICV_4 $T=73140 198560 1 0 $X=72950 $Y=195600
X490 1 2 405 ICV_4 $T=73140 214880 1 0 $X=72950 $Y=211920
X491 1 2 80 ICV_4 $T=90160 187680 1 0 $X=89970 $Y=184720
X492 1 2 73 ICV_4 $T=94300 204000 0 0 $X=94110 $Y=203760
X493 1 2 82 ICV_4 $T=98900 204000 1 0 $X=98710 $Y=201040
X494 1 2 419 ICV_4 $T=113160 193120 0 0 $X=112970 $Y=192880
X495 1 2 427 ICV_4 $T=114540 198560 0 0 $X=114350 $Y=198320
X496 1 2 99 ICV_4 $T=123740 176800 1 0 $X=123550 $Y=173840
X497 1 2 435 ICV_4 $T=124660 198560 0 0 $X=124470 $Y=198320
X498 1 2 104 ICV_4 $T=131560 187680 0 0 $X=131370 $Y=187440
X499 1 2 99 ICV_4 $T=132940 176800 0 0 $X=132750 $Y=176560
X500 1 2 90 ICV_4 $T=133400 214880 1 0 $X=133210 $Y=211920
X501 1 2 436 ICV_4 $T=134320 204000 1 0 $X=134130 $Y=201040
X502 1 2 106 ICV_4 $T=134320 209440 1 0 $X=134130 $Y=206480
X503 1 2 110 ICV_4 $T=141220 214880 0 0 $X=141030 $Y=214640
X504 1 2 114 ICV_4 $T=143060 176800 0 0 $X=142870 $Y=176560
X505 1 2 97 ICV_4 $T=147200 214880 0 0 $X=147010 $Y=214640
X506 1 2 448 ICV_4 $T=148580 209440 1 0 $X=148390 $Y=206480
X507 1 2 102 ICV_4 $T=152720 176800 0 0 $X=152530 $Y=176560
X508 1 2 466 ICV_4 $T=179860 204000 1 0 $X=179670 $Y=201040
X509 1 2 153 ICV_4 $T=192280 187680 0 0 $X=192090 $Y=187440
X510 1 2 159 ICV_4 $T=195040 193120 0 0 $X=194850 $Y=192880
X511 1 2 163 ICV_4 $T=198720 176800 0 0 $X=198530 $Y=176560
X512 1 2 471 ICV_4 $T=205160 198560 1 0 $X=204970 $Y=195600
X513 1 2 182 ICV_4 $T=217580 204000 0 0 $X=217390 $Y=203760
X514 1 2 186 ICV_4 $T=217580 209440 0 0 $X=217390 $Y=209200
X515 1 2 190 ICV_4 $T=223560 182240 1 0 $X=223370 $Y=179280
X516 1 2 182 ICV_4 $T=227240 204000 0 0 $X=227050 $Y=203760
X517 1 2 196 ICV_4 $T=237360 176800 1 0 $X=237170 $Y=173840
X518 1 2 200 ICV_4 $T=237360 182240 1 0 $X=237170 $Y=179280
X519 1 2 4 ICV_4 $T=245640 182240 0 0 $X=245450 $Y=182000
X520 1 2 495 ICV_4 $T=249320 182240 1 0 $X=249130 $Y=179280
X521 1 2 203 ICV_4 $T=254840 209440 0 0 $X=254650 $Y=209200
X522 1 2 207 ICV_4 $T=256220 209440 1 0 $X=256030 $Y=206480
X523 1 2 229 ICV_4 $T=278760 214880 1 0 $X=278570 $Y=211920
X524 1 2 229 ICV_4 $T=281980 214880 1 0 $X=281790 $Y=211920
X525 1 2 510 ICV_4 $T=283360 187680 0 0 $X=283170 $Y=187440
X526 1 2 505 ICV_4 $T=283360 193120 0 0 $X=283170 $Y=192880
X527 1 2 231 ICV_4 $T=283360 214880 0 0 $X=283170 $Y=214640
X528 1 2 232 ICV_4 $T=284740 209440 1 0 $X=284550 $Y=206480
X529 1 2 4 ICV_4 $T=287500 209440 1 0 $X=287310 $Y=206480
X530 1 2 514 ICV_4 $T=289340 176800 0 0 $X=289150 $Y=176560
X531 1 2 518 ICV_4 $T=297620 187680 1 0 $X=297430 $Y=184720
X532 1 2 521 ICV_4 $T=298080 176800 0 0 $X=297890 $Y=176560
X533 1 2 222 ICV_4 $T=299000 209440 0 0 $X=298810 $Y=209200
X534 1 2 250 ICV_4 $T=304980 214880 1 0 $X=304790 $Y=211920
X535 1 2 439 ICV_4 $T=309120 187680 0 0 $X=308930 $Y=187440
X536 1 2 523 ICV_4 $T=310500 209440 1 0 $X=310310 $Y=206480
X537 1 2 4 ICV_4 $T=311420 214880 0 0 $X=311230 $Y=214640
X538 1 2 248 ICV_4 $T=317860 214880 1 0 $X=317670 $Y=211920
X539 1 2 426 ICV_4 $T=339480 198560 0 0 $X=339290 $Y=198320
X540 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 182240 1 0 $X=16370 $Y=179280
X541 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=18400 214880 0 0 $X=18210 $Y=214640
X542 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=28980 176800 0 0 $X=28790 $Y=176560
X543 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30820 182240 1 0 $X=30630 $Y=179280
X544 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=30820 204000 0 0 $X=30630 $Y=203760
X545 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=33120 187680 1 0 $X=32930 $Y=184720
X546 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 176800 1 0 $X=48110 $Y=173840
X547 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=51520 198560 0 0 $X=51330 $Y=198320
X548 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=53820 204000 1 0 $X=53630 $Y=201040
X549 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=59340 182240 1 0 $X=59150 $Y=179280
X550 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 204000 1 0 $X=72490 $Y=201040
X551 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=81420 198560 0 0 $X=81230 $Y=198320
X552 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 182240 0 0 $X=89970 $Y=182000
X553 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 214880 0 0 $X=89970 $Y=214640
X554 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=92460 214880 1 0 $X=92270 $Y=211920
X555 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101200 209440 1 0 $X=101010 $Y=206480
X556 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101660 176800 0 0 $X=101470 $Y=176560
X557 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=109480 204000 1 0 $X=109290 $Y=201040
X558 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=112700 182240 0 0 $X=112510 $Y=182000
X559 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=120980 193120 1 0 $X=120790 $Y=190160
X560 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=127420 214880 1 0 $X=127230 $Y=211920
X561 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=142600 198560 0 0 $X=142410 $Y=198320
X562 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 187680 0 0 $X=142870 $Y=187440
X563 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=145360 193120 1 0 $X=145170 $Y=190160
X564 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157320 182240 1 0 $X=157130 $Y=179280
X565 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=164220 214880 0 0 $X=164030 $Y=214640
X566 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=165140 176800 0 0 $X=164950 $Y=176560
X567 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=168360 176800 1 0 $X=168170 $Y=173840
X568 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=168820 198560 0 0 $X=168630 $Y=198320
X569 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=172040 204000 1 0 $X=171850 $Y=201040
X570 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=172500 214880 1 0 $X=172310 $Y=211920
X571 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=184920 187680 1 0 $X=184730 $Y=184720
X572 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 193120 0 0 $X=185190 $Y=192880
X573 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=186300 214880 0 0 $X=186110 $Y=214640
X574 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=188600 209440 1 0 $X=188410 $Y=206480
X575 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=195040 176800 1 0 $X=194850 $Y=173840
X576 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=198720 182240 0 0 $X=198530 $Y=182000
X577 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=204240 214880 1 0 $X=204050 $Y=211920
X578 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=227700 193120 1 0 $X=227510 $Y=190160
X579 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=247480 193120 0 0 $X=247290 $Y=192880
X580 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=247480 198560 1 0 $X=247290 $Y=195600
X581 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=253460 193120 0 0 $X=253270 $Y=192880
X582 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=255760 193120 1 0 $X=255570 $Y=190160
X583 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=267260 187680 1 0 $X=267070 $Y=184720
X584 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=285200 204000 1 0 $X=285010 $Y=201040
X585 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=286580 176800 0 0 $X=286390 $Y=176560
X586 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=311420 187680 1 0 $X=311230 $Y=184720
X587 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331200 182240 0 0 $X=331010 $Y=182000
X588 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331660 187680 0 0 $X=331470 $Y=187440
X589 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339020 204000 0 0 $X=338830 $Y=203760
X590 1 2 33 ICV_5 $T=43700 187680 0 0 $X=43510 $Y=187440
X591 1 2 52 ICV_5 $T=65320 176800 0 0 $X=65130 $Y=176560
X592 1 2 407 ICV_5 $T=77280 198560 1 0 $X=77090 $Y=195600
X593 1 2 70 ICV_5 $T=79580 209440 0 0 $X=79390 $Y=209200
X594 1 2 411 ICV_5 $T=84180 193120 0 0 $X=83990 $Y=192880
X595 1 2 40 ICV_5 $T=86020 182240 0 0 $X=85830 $Y=182000
X596 1 2 86 ICV_5 $T=105340 176800 1 0 $X=105150 $Y=173840
X597 1 2 371 ICV_5 $T=127880 198560 1 0 $X=127690 $Y=195600
X598 1 2 453 ICV_5 $T=166060 193120 1 0 $X=165870 $Y=190160
X599 1 2 131 ICV_5 $T=168360 176800 0 0 $X=168170 $Y=176560
X600 1 2 49 ICV_5 $T=220800 209440 0 0 $X=220610 $Y=209200
X601 1 2 4 ICV_5 $T=230460 193120 1 0 $X=230270 $Y=190160
X602 1 2 482 ICV_5 $T=230920 204000 1 0 $X=230730 $Y=201040
X603 1 2 485 ICV_5 $T=235060 204000 0 0 $X=234870 $Y=203760
X604 1 2 172 ICV_5 $T=237820 209440 0 0 $X=237630 $Y=209200
X605 1 2 174 ICV_5 $T=240120 182240 1 0 $X=239930 $Y=179280
X606 1 2 489 ICV_5 $T=240120 204000 1 0 $X=239930 $Y=201040
X607 1 2 201 ICV_5 $T=240580 176800 1 0 $X=240390 $Y=173840
X608 1 2 120 ICV_5 $T=282440 176800 0 0 $X=282250 $Y=176560
X609 1 2 372 ICV_5 $T=320620 193120 0 0 $X=320430 $Y=192880
X610 1 2 532 ICV_5 $T=324760 209440 1 0 $X=324570 $Y=206480
X611 1 2 449 ICV_5 $T=338100 187680 0 0 $X=337910 $Y=187440
X612 1 2 3 ICV_5 $T=338100 214880 0 0 $X=337910 $Y=214640
X613 1 2 20 ICV_6 $T=40480 204000 1 0 $X=40290 $Y=201040
X614 1 2 397 ICV_6 $T=49220 209440 1 0 $X=49030 $Y=206480
X615 1 2 44 ICV_6 $T=51980 209440 0 0 $X=51790 $Y=209200
X616 1 2 406 ICV_6 $T=68080 193120 1 0 $X=67890 $Y=190160
X617 1 2 62 ICV_6 $T=69920 209440 1 0 $X=69730 $Y=206480
X618 1 2 408 ICV_6 $T=71300 182240 1 0 $X=71110 $Y=179280
X619 1 2 407 ICV_6 $T=80960 187680 0 0 $X=80770 $Y=187440
X620 1 2 42 ICV_6 $T=91080 176800 0 0 $X=90890 $Y=176560
X621 1 2 79 ICV_6 $T=92920 182240 0 0 $X=92730 $Y=182000
X622 1 2 413 ICV_6 $T=97980 187680 1 0 $X=97790 $Y=184720
X623 1 2 430 ICV_6 $T=118220 182240 1 0 $X=118030 $Y=179280
X624 1 2 100 ICV_6 $T=123740 214880 0 0 $X=123550 $Y=214640
X625 1 2 113 ICV_6 $T=138460 182240 1 0 $X=138270 $Y=179280
X626 1 2 4 ICV_6 $T=140760 204000 0 0 $X=140570 $Y=203760
X627 1 2 127 ICV_6 $T=155480 176800 1 0 $X=155290 $Y=173840
X628 1 2 449 ICV_6 $T=165600 182240 0 0 $X=165410 $Y=182000
X629 1 2 454 ICV_6 $T=166060 198560 1 0 $X=165870 $Y=195600
X630 1 2 136 ICV_6 $T=177560 209440 1 0 $X=177370 $Y=206480
X631 1 2 144 ICV_6 $T=187680 209440 0 0 $X=187490 $Y=209200
X632 1 2 81 ICV_6 $T=194580 198560 0 0 $X=194390 $Y=198320
X633 1 2 69 ICV_6 $T=195040 187680 0 0 $X=194850 $Y=187440
X634 1 2 181 ICV_6 $T=210680 176800 1 0 $X=210490 $Y=173840
X635 1 2 484 ICV_6 $T=230460 214880 1 0 $X=230270 $Y=211920
X636 1 2 502 ICV_6 $T=266800 182240 1 0 $X=266610 $Y=179280
X637 1 2 218 ICV_6 $T=267720 209440 1 0 $X=267530 $Y=206480
X638 1 2 225 ICV_6 $T=275080 176800 0 0 $X=274890 $Y=176560
X639 1 2 517 ICV_6 $T=294400 198560 1 0 $X=294210 $Y=195600
X640 1 2 240 ICV_6 $T=294400 204000 1 0 $X=294210 $Y=201040
X641 1 2 520 ICV_6 $T=304520 176800 0 0 $X=304330 $Y=176560
X642 1 2 242 ICV_6 $T=304520 209440 1 0 $X=304330 $Y=206480
X643 1 2 262 ICV_6 $T=337640 176800 0 0 $X=337450 $Y=176560
X644 1 2 530 ICV_6 $T=337640 182240 0 0 $X=337450 $Y=182000
X645 1 2 495 ICV_6 $T=343620 193120 0 0 $X=343430 $Y=192880
X646 1 3 5 ICV_7 $T=7820 176800 1 0 $X=7630 $Y=173840
X647 1 3 4 ICV_7 $T=7820 187680 1 0 $X=7630 $Y=184720
X648 1 3 4 ICV_7 $T=7820 193120 1 0 $X=7630 $Y=190160
X649 1 3 373 ICV_7 $T=7820 198560 1 0 $X=7630 $Y=195600
X650 1 3 4 ICV_7 $T=7820 209440 1 0 $X=7630 $Y=206480
X651 1 3 4 ICV_7 $T=7820 214880 1 0 $X=7630 $Y=211920
X652 1 377 16 ICV_7 $T=21160 209440 1 0 $X=20970 $Y=206480
X653 1 17 20 ICV_7 $T=23460 193120 1 0 $X=23270 $Y=190160
X654 1 378 15 ICV_7 $T=26220 176800 0 0 $X=26030 $Y=176560
X655 1 380 385 ICV_7 $T=26220 198560 0 0 $X=26030 $Y=198320
X656 1 383 16 ICV_7 $T=27140 182240 0 0 $X=26950 $Y=182000
X657 1 4 384 ICV_7 $T=27140 187680 0 0 $X=26950 $Y=187440
X658 1 386 23 ICV_7 $T=28060 209440 0 0 $X=27870 $Y=209200
X659 1 387 14 ICV_7 $T=29900 198560 0 0 $X=29710 $Y=198320
X660 1 24 26 ICV_7 $T=29900 214880 0 0 $X=29710 $Y=214640
X661 1 380 23 ICV_7 $T=34960 187680 0 0 $X=34770 $Y=187440
X662 1 17 394 ICV_7 $T=36800 204000 1 0 $X=36610 $Y=201040
X663 1 28 388 ICV_7 $T=38640 176800 1 0 $X=38450 $Y=173840
X664 1 395 395 ICV_7 $T=43700 193120 1 0 $X=43510 $Y=190160
X665 1 390 23 ICV_7 $T=48300 209440 0 0 $X=48110 $Y=209200
X666 1 42 40 ICV_7 $T=48760 182240 0 0 $X=48570 $Y=182000
X667 1 396 390 ICV_7 $T=50140 193120 0 0 $X=49950 $Y=192880
X668 1 399 400 ICV_7 $T=50600 198560 1 0 $X=50410 $Y=195600
X669 1 398 45 ICV_7 $T=51980 214880 0 0 $X=51790 $Y=214640
X670 1 4 402 ICV_7 $T=55200 182240 0 0 $X=55010 $Y=182000
X671 1 47 44 ICV_7 $T=55200 204000 0 0 $X=55010 $Y=203760
X672 1 53 57 ICV_7 $T=63020 214880 1 0 $X=62830 $Y=211920
X673 1 55 396 ICV_7 $T=64400 193120 1 0 $X=64210 $Y=190160
X674 1 26 4 ICV_7 $T=64400 209440 0 0 $X=64210 $Y=209200
X675 1 405 61 ICV_7 $T=66240 209440 1 0 $X=66050 $Y=206480
X676 1 33 56 ICV_7 $T=68080 187680 0 0 $X=67890 $Y=187440
X677 1 67 50 ICV_7 $T=76360 204000 0 0 $X=76170 $Y=203760
X678 1 69 404 ICV_7 $T=77280 187680 0 0 $X=77090 $Y=187440
X679 1 4 71 ICV_7 $T=77740 214880 0 0 $X=77550 $Y=214640
X680 1 409 73 ICV_7 $T=80500 193120 0 0 $X=80310 $Y=192880
X681 1 412 64 ICV_7 $T=84180 198560 0 0 $X=83990 $Y=198320
X682 1 413 78 ICV_7 $T=86020 187680 0 0 $X=85830 $Y=187440
X683 1 76 415 ICV_7 $T=86020 204000 0 0 $X=85830 $Y=203760
X684 1 414 65 ICV_7 $T=87400 198560 1 0 $X=87210 $Y=195600
X685 1 64 419 ICV_7 $T=91080 193120 0 0 $X=90890 $Y=192880
X686 1 82 78 ICV_7 $T=97520 193120 1 0 $X=97330 $Y=190160
X687 1 420 425 ICV_7 $T=98440 198560 1 0 $X=98250 $Y=195600
X688 1 423 425 ICV_7 $T=98440 209440 1 0 $X=98250 $Y=206480
X689 1 84 50 ICV_7 $T=98900 176800 0 0 $X=98710 $Y=176560
X690 1 81 404 ICV_7 $T=105340 193120 1 0 $X=105150 $Y=190160
X691 1 90 4 ICV_7 $T=110860 198560 0 0 $X=110670 $Y=198320
X692 1 428 90 ICV_7 $T=114080 204000 0 0 $X=113890 $Y=203760
X693 1 431 33 ICV_7 $T=120060 176800 0 0 $X=119870 $Y=176560
X694 1 95 96 ICV_7 $T=120060 214880 0 0 $X=119870 $Y=214640
X695 1 95 95 ICV_7 $T=120520 204000 0 0 $X=120330 $Y=203760
X696 1 433 434 ICV_7 $T=124200 204000 1 0 $X=124010 $Y=201040
X697 1 433 101 ICV_7 $T=124660 214880 1 0 $X=124470 $Y=211920
X698 1 436 94 ICV_7 $T=127880 204000 1 0 $X=127690 $Y=201040
X699 1 437 108 ICV_7 $T=128340 214880 0 0 $X=128150 $Y=214640
X700 1 105 109 ICV_7 $T=129260 176800 0 0 $X=129070 $Y=176560
X701 1 110 111 ICV_7 $T=131100 209440 0 0 $X=130910 $Y=209200
X702 1 4 440 ICV_7 $T=134780 187680 0 0 $X=134590 $Y=187440
X703 1 116 118 ICV_7 $T=141220 214880 1 0 $X=141030 $Y=211920
X704 1 445 4 ICV_7 $T=146740 187680 1 0 $X=146550 $Y=184720
X705 1 443 94 ICV_7 $T=154560 209440 0 0 $X=154370 $Y=209200
X706 1 4 451 ICV_7 $T=160540 198560 0 0 $X=160350 $Y=198320
X707 1 4 452 ICV_7 $T=161920 209440 0 0 $X=161730 $Y=209200
X708 1 132 4 ICV_7 $T=167440 214880 0 0 $X=167250 $Y=214640
X709 1 455 460 ICV_7 $T=169740 193120 1 0 $X=169550 $Y=190160
X710 1 456 459 ICV_7 $T=170200 182240 0 0 $X=170010 $Y=182000
X711 1 457 137 ICV_7 $T=170200 204000 0 0 $X=170010 $Y=203760
X712 1 458 460 ICV_7 $T=170660 198560 1 0 $X=170470 $Y=195600
X713 1 463 4 ICV_7 $T=174340 176800 1 0 $X=174150 $Y=173840
X714 1 139 140 ICV_7 $T=175260 198560 0 0 $X=175070 $Y=198320
X715 1 142 139 ICV_7 $T=181700 187680 0 0 $X=181510 $Y=187440
X716 1 139 465 ICV_7 $T=182160 187680 1 0 $X=181970 $Y=184720
X717 1 130 462 ICV_7 $T=182620 176800 0 0 $X=182430 $Y=176560
X718 1 462 466 ICV_7 $T=182620 193120 0 0 $X=182430 $Y=192880
X719 1 152 148 ICV_7 $T=189520 214880 0 0 $X=189330 $Y=214640
X720 1 4 160 ICV_7 $T=193660 209440 0 0 $X=193470 $Y=209200
X721 1 166 4 ICV_7 $T=198260 193120 0 0 $X=198070 $Y=192880
X722 1 167 168 ICV_7 $T=198260 214880 0 0 $X=198070 $Y=214640
X723 1 174 470 ICV_7 $T=203320 187680 0 0 $X=203130 $Y=187440
X724 1 469 52 ICV_7 $T=203780 182240 1 0 $X=203590 $Y=179280
X725 1 177 48 ICV_7 $T=207000 214880 1 0 $X=206810 $Y=211920
X726 1 50 472 ICV_7 $T=207460 182240 1 0 $X=207270 $Y=179280
X727 1 178 473 ICV_7 $T=208380 198560 1 0 $X=208190 $Y=195600
X728 1 182 177 ICV_7 $T=210680 214880 1 0 $X=210490 $Y=211920
X729 1 184 474 ICV_7 $T=213900 209440 0 0 $X=213710 $Y=209200
X730 1 171 477 ICV_7 $T=216660 198560 0 0 $X=216470 $Y=198320
X731 1 183 480 ICV_7 $T=219880 204000 1 0 $X=219690 $Y=201040
X732 1 478 182 ICV_7 $T=221720 198560 1 0 $X=221530 $Y=195600
X733 1 189 182 ICV_7 $T=221720 214880 0 0 $X=221530 $Y=214640
X734 1 479 174 ICV_7 $T=222180 176800 0 0 $X=221990 $Y=176560
X735 1 481 483 ICV_7 $T=224480 193120 0 0 $X=224290 $Y=192880
X736 1 122 194 ICV_7 $T=224480 209440 0 0 $X=224290 $Y=209200
X737 1 183 480 ICV_7 $T=225400 198560 1 0 $X=225210 $Y=195600
X738 1 192 191 ICV_7 $T=226320 176800 0 0 $X=226130 $Y=176560
X739 1 183 484 ICV_7 $T=231380 204000 0 0 $X=231190 $Y=203760
X740 1 486 197 ICV_7 $T=233680 176800 0 0 $X=233490 $Y=176560
X741 1 199 4 ICV_7 $T=236440 198560 0 0 $X=236250 $Y=198320
X742 1 488 202 ICV_7 $T=239200 204000 0 0 $X=239010 $Y=203760
X743 1 54 493 ICV_7 $T=241500 209440 0 0 $X=241310 $Y=209200
X744 1 490 207 ICV_7 $T=245180 214880 0 0 $X=244990 $Y=214640
X745 1 492 206 ICV_7 $T=245640 182240 1 0 $X=245450 $Y=179280
X746 1 202 496 ICV_7 $T=250700 193120 0 0 $X=250510 $Y=192880
X747 1 494 171 ICV_7 $T=251620 204000 1 0 $X=251430 $Y=201040
X748 1 4 497 ICV_7 $T=252540 176800 0 0 $X=252350 $Y=176560
X749 1 498 216 ICV_7 $T=258520 193120 1 0 $X=258330 $Y=190160
X750 1 4 500 ICV_7 $T=259440 198560 0 0 $X=259250 $Y=198320
X751 1 202 499 ICV_7 $T=259440 204000 0 0 $X=259250 $Y=203760
X752 1 213 210 ICV_7 $T=259440 214880 0 0 $X=259250 $Y=214640
X753 1 172 4 ICV_7 $T=264040 209440 0 0 $X=263850 $Y=209200
X754 1 501 439 ICV_7 $T=265420 187680 0 0 $X=265230 $Y=187440
X755 1 220 4 ICV_7 $T=270940 193120 0 0 $X=270750 $Y=192880
X756 1 439 506 ICV_7 $T=273700 198560 0 0 $X=273510 $Y=198320
X757 1 120 510 ICV_7 $T=278300 182240 0 0 $X=278110 $Y=182000
X758 1 509 507 ICV_7 $T=281980 182240 0 0 $X=281790 $Y=182000
X759 1 222 511 ICV_7 $T=282440 209440 0 0 $X=282250 $Y=209200
X760 1 146 234 ICV_7 $T=287960 198560 0 0 $X=287770 $Y=198320
X761 1 513 509 ICV_7 $T=288420 182240 1 0 $X=288230 $Y=179280
X762 1 220 515 ICV_7 $T=288420 193120 1 0 $X=288230 $Y=190160
X763 1 512 510 ICV_7 $T=290720 193120 0 0 $X=290530 $Y=192880
X764 1 239 237 ICV_7 $T=294400 176800 0 0 $X=294210 $Y=176560
X765 1 510 510 ICV_7 $T=294400 182240 0 0 $X=294210 $Y=182000
X766 1 238 509 ICV_7 $T=294400 193120 1 0 $X=294210 $Y=190160
X767 1 520 509 ICV_7 $T=296240 182240 1 0 $X=296050 $Y=179280
X768 1 164 220 ICV_7 $T=300840 176800 0 0 $X=300650 $Y=176560
X769 1 243 249 ICV_7 $T=301300 214880 0 0 $X=301110 $Y=214640
X770 1 439 522 ICV_7 $T=305440 182240 0 0 $X=305250 $Y=182000
X771 1 244 249 ICV_7 $T=306820 209440 0 0 $X=306630 $Y=209200
X772 1 252 526 ICV_7 $T=307740 198560 0 0 $X=307550 $Y=198320
X773 1 524 4 ICV_7 $T=310500 176800 0 0 $X=310310 $Y=176560
X774 1 4 527 ICV_7 $T=310500 193120 0 0 $X=310310 $Y=192880
X775 1 248 246 ICV_7 $T=310500 209440 0 0 $X=310310 $Y=209200
X776 1 525 530 ICV_7 $T=314640 187680 1 0 $X=314450 $Y=184720
X777 1 250 528 ICV_7 $T=315560 198560 0 0 $X=315370 $Y=198320
X778 1 248 246 ICV_7 $T=315560 204000 0 0 $X=315370 $Y=203760
X779 1 252 531 ICV_7 $T=321080 209440 1 0 $X=320890 $Y=206480
X780 1 533 260 ICV_7 $T=322000 198560 1 0 $X=321810 $Y=195600
X781 1 246 533 ICV_7 $T=322000 204000 1 0 $X=321810 $Y=201040
X782 1 3 4 ICV_7 $T=333960 176800 0 0 $X=333770 $Y=176560
X783 1 3 4 ICV_7 $T=333960 182240 0 0 $X=333770 $Y=182000
X784 1 3 4 ICV_7 $T=334420 187680 0 0 $X=334230 $Y=187440
X785 1 4 263 ICV_7 $T=334880 214880 1 0 $X=334690 $Y=211920
X786 1 3 4 ICV_7 $T=335800 198560 0 0 $X=335610 $Y=198320
X787 1 2 3 5 4 2 7 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 176800 0 0 $X=7630 $Y=176560
X788 1 2 3 371 4 2 8 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 187680 0 0 $X=7630 $Y=187440
X789 1 2 3 372 4 2 9 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 193120 0 0 $X=7630 $Y=192880
X790 1 2 3 373 4 2 10 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 198560 0 0 $X=7630 $Y=198320
X791 1 2 3 370 4 2 11 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 209440 0 0 $X=7630 $Y=209200
X792 1 2 3 6 4 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 214880 0 0 $X=7630 $Y=214640
X793 1 2 537 374 4 2 15 1 sky130_fd_sc_hd__dfrtp_4 $T=10120 182240 0 0 $X=9930 $Y=182000
X794 1 2 538 376 4 2 373 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 198560 1 0 $X=20970 $Y=195600
X795 1 2 539 377 4 2 370 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 214880 1 0 $X=20970 $Y=211920
X796 1 2 540 384 4 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=27140 193120 1 0 $X=26950 $Y=190160
X797 1 2 541 393 4 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=33580 209440 1 0 $X=33390 $Y=206480
X798 1 2 542 402 4 2 56 1 sky130_fd_sc_hd__dfrtp_4 $T=55200 187680 1 0 $X=55010 $Y=184720
X799 1 2 543 403 4 2 58 1 sky130_fd_sc_hd__dfrtp_4 $T=56580 204000 1 0 $X=56390 $Y=201040
X800 1 2 544 61 4 2 70 1 sky130_fd_sc_hd__dfrtp_4 $T=68080 209440 0 0 $X=67890 $Y=209200
X801 1 2 545 408 4 2 72 1 sky130_fd_sc_hd__dfrtp_4 $T=71300 176800 0 0 $X=71110 $Y=176560
X802 1 2 546 410 4 2 79 1 sky130_fd_sc_hd__dfrtp_4 $T=78660 187680 1 0 $X=78470 $Y=184720
X803 1 2 547 421 4 2 85 1 sky130_fd_sc_hd__dfrtp_4 $T=95220 214880 0 0 $X=95030 $Y=214640
X804 1 2 548 420 4 2 426 1 sky130_fd_sc_hd__dfrtp_4 $T=98440 198560 0 0 $X=98250 $Y=198320
X805 1 2 549 423 4 2 88 1 sky130_fd_sc_hd__dfrtp_4 $T=98440 209440 0 0 $X=98250 $Y=209200
X806 1 2 550 87 4 2 89 1 sky130_fd_sc_hd__dfrtp_4 $T=105340 182240 1 0 $X=105150 $Y=179280
X807 1 2 551 427 4 2 371 1 sky130_fd_sc_hd__dfrtp_4 $T=112700 204000 1 0 $X=112510 $Y=201040
X808 1 2 552 429 4 2 98 1 sky130_fd_sc_hd__dfrtp_4 $T=116380 198560 1 0 $X=116190 $Y=195600
X809 1 2 553 430 4 2 103 1 sky130_fd_sc_hd__dfrtp_4 $T=119140 182240 0 0 $X=118950 $Y=182000
X810 1 2 554 440 4 2 117 1 sky130_fd_sc_hd__dfrtp_4 $T=134780 193120 1 0 $X=134590 $Y=190160
X811 1 2 555 441 4 2 121 1 sky130_fd_sc_hd__dfrtp_4 $T=137080 209440 1 0 $X=136890 $Y=206480
X812 1 2 556 445 4 2 127 1 sky130_fd_sc_hd__dfrtp_4 $T=147200 182240 0 0 $X=147010 $Y=182000
X813 1 2 557 448 4 2 126 1 sky130_fd_sc_hd__dfrtp_4 $T=148120 204000 0 0 $X=147930 $Y=203760
X814 1 2 558 447 4 2 449 1 sky130_fd_sc_hd__dfrtp_4 $T=148580 187680 0 0 $X=148390 $Y=187440
X815 1 2 559 450 4 2 131 1 sky130_fd_sc_hd__dfrtp_4 $T=161460 187680 1 0 $X=161270 $Y=184720
X816 1 2 560 451 4 2 133 1 sky130_fd_sc_hd__dfrtp_4 $T=161460 204000 1 0 $X=161270 $Y=201040
X817 1 2 561 452 4 2 136 1 sky130_fd_sc_hd__dfrtp_4 $T=161920 214880 1 0 $X=161730 $Y=211920
X818 1 2 562 138 4 2 147 1 sky130_fd_sc_hd__dfrtp_4 $T=175720 214880 0 0 $X=175530 $Y=214640
X819 1 2 563 160 4 2 167 1 sky130_fd_sc_hd__dfrtp_4 $T=193660 214880 1 0 $X=193470 $Y=211920
X820 1 2 564 468 4 2 170 1 sky130_fd_sc_hd__dfrtp_4 $T=203320 193120 0 0 $X=203130 $Y=192880
X821 1 2 565 471 4 2 179 1 sky130_fd_sc_hd__dfrtp_4 $T=205160 198560 0 0 $X=204970 $Y=198320
X822 1 2 566 181 4 2 188 1 sky130_fd_sc_hd__dfrtp_4 $T=210680 176800 0 0 $X=210490 $Y=176560
X823 1 2 567 476 4 2 190 1 sky130_fd_sc_hd__dfrtp_4 $T=217580 187680 1 0 $X=217390 $Y=184720
X824 1 2 568 481 4 2 199 1 sky130_fd_sc_hd__dfrtp_4 $T=229080 198560 1 0 $X=228890 $Y=195600
X825 1 2 569 483 4 2 198 1 sky130_fd_sc_hd__dfrtp_4 $T=231380 193120 0 0 $X=231190 $Y=192880
X826 1 2 570 489 4 2 205 1 sky130_fd_sc_hd__dfrtp_4 $T=240120 198560 0 0 $X=239930 $Y=198320
X827 1 2 571 492 4 2 495 1 sky130_fd_sc_hd__dfrtp_4 $T=245640 187680 1 0 $X=245450 $Y=184720
X828 1 2 572 497 4 2 212 1 sky130_fd_sc_hd__dfrtp_4 $T=252080 182240 1 0 $X=251890 $Y=179280
X829 1 2 573 500 4 2 217 1 sky130_fd_sc_hd__dfrtp_4 $T=258060 204000 1 0 $X=257870 $Y=201040
X830 1 2 574 498 4 2 216 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 193120 0 0 $X=259250 $Y=192880
X831 1 2 575 502 4 2 225 1 sky130_fd_sc_hd__dfrtp_4 $T=266800 182240 0 0 $X=266610 $Y=182000
X832 1 2 576 218 4 2 223 1 sky130_fd_sc_hd__dfrtp_4 $T=267720 209440 0 0 $X=267530 $Y=209200
X833 1 2 577 504 4 2 228 1 sky130_fd_sc_hd__dfrtp_4 $T=273700 198560 1 0 $X=273510 $Y=195600
X834 1 2 578 511 4 2 240 1 sky130_fd_sc_hd__dfrtp_4 $T=287500 209440 0 0 $X=287310 $Y=209200
X835 1 2 579 516 4 2 242 1 sky130_fd_sc_hd__dfrtp_4 $T=290720 204000 0 0 $X=290530 $Y=203760
X836 1 2 580 518 4 2 247 1 sky130_fd_sc_hd__dfrtp_4 $T=297620 187680 0 0 $X=297430 $Y=187440
X837 1 2 581 254 4 2 251 1 sky130_fd_sc_hd__dfrtp_4 $T=308200 176800 1 0 $X=308010 $Y=173840
X838 1 2 582 527 4 2 372 1 sky130_fd_sc_hd__dfrtp_4 $T=310500 198560 1 0 $X=310310 $Y=195600
X839 1 2 583 524 4 2 257 1 sky130_fd_sc_hd__dfrtp_4 $T=315560 176800 0 0 $X=315370 $Y=176560
X840 1 2 584 525 4 2 530 1 sky130_fd_sc_hd__dfrtp_4 $T=315560 187680 0 0 $X=315370 $Y=187440
X841 1 2 585 535 4 2 261 1 sky130_fd_sc_hd__dfrtp_4 $T=326140 193120 0 0 $X=325950 $Y=192880
X842 1 2 586 536 4 2 263 1 sky130_fd_sc_hd__dfrtp_4 $T=326600 214880 0 0 $X=326410 $Y=214640
X843 1 2 3 216 4 2 264 1 sky130_fd_sc_hd__dfrtp_4 $T=333960 176800 1 0 $X=333770 $Y=173840
X844 1 2 3 262 4 2 265 1 sky130_fd_sc_hd__dfrtp_4 $T=333960 182240 1 0 $X=333770 $Y=179280
X845 1 2 3 530 4 2 266 1 sky130_fd_sc_hd__dfrtp_4 $T=333960 187680 1 0 $X=333770 $Y=184720
X846 1 2 3 449 4 2 267 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 193120 1 0 $X=334230 $Y=190160
X847 1 2 3 495 4 2 268 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 198560 1 0 $X=334690 $Y=195600
X848 1 2 3 426 4 2 269 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 204000 1 0 $X=334690 $Y=201040
X849 1 2 388 ICV_13 $T=29900 182240 0 0 $X=29710 $Y=182000
X850 1 2 389 ICV_13 $T=29900 187680 0 0 $X=29710 $Y=187440
X851 1 2 25 ICV_13 $T=29900 193120 0 0 $X=29710 $Y=192880
X852 1 2 38 ICV_13 $T=41400 176800 1 0 $X=41210 $Y=173840
X853 1 2 39 ICV_13 $T=42320 198560 0 0 $X=42130 $Y=198320
X854 1 2 404 ICV_13 $T=57960 193120 0 0 $X=57770 $Y=192880
X855 1 2 81 ICV_13 $T=90160 187680 0 0 $X=89970 $Y=187440
X856 1 2 414 ICV_13 $T=100280 193120 1 0 $X=100090 $Y=190160
X857 1 2 83 ICV_13 $T=103040 193120 0 0 $X=102850 $Y=192880
X858 1 2 97 ICV_13 $T=120980 209440 0 0 $X=120790 $Y=209200
X859 1 2 438 ICV_13 $T=128340 176800 1 0 $X=128150 $Y=173840
X860 1 2 107 ICV_13 $T=128340 209440 1 0 $X=128150 $Y=206480
X861 1 2 97 ICV_13 $T=130640 204000 0 0 $X=130450 $Y=203760
X862 1 2 95 ICV_13 $T=142140 209440 0 0 $X=141950 $Y=209200
X863 1 2 135 ICV_13 $T=170200 187680 0 0 $X=170010 $Y=187440
X864 1 2 462 ICV_13 $T=170200 193120 0 0 $X=170010 $Y=192880
X865 1 2 138 ICV_13 $T=170200 214880 0 0 $X=170010 $Y=214640
X866 1 2 460 ICV_13 $T=184460 176800 1 0 $X=184270 $Y=173840
X867 1 2 149 ICV_13 $T=184460 182240 1 0 $X=184270 $Y=179280
X868 1 2 158 ICV_13 $T=192740 176800 0 0 $X=192550 $Y=176560
X869 1 2 474 ICV_13 $T=212520 204000 1 0 $X=212330 $Y=201040
X870 1 2 178 ICV_13 $T=226320 198560 0 0 $X=226130 $Y=198320
X871 1 2 204 ICV_13 $T=243800 176800 0 0 $X=243610 $Y=176560
X872 1 2 205 ICV_13 $T=244720 198560 1 0 $X=244530 $Y=195600
X873 1 2 203 ICV_13 $T=247020 204000 0 0 $X=246830 $Y=203760
X874 1 2 211 ICV_13 $T=254380 214880 0 0 $X=254190 $Y=214640
X875 1 2 162 ICV_13 $T=273240 187680 0 0 $X=273050 $Y=187440
X876 1 2 509 ICV_13 $T=275080 187680 1 0 $X=274890 $Y=184720
X877 1 2 236 ICV_13 $T=288880 214880 1 0 $X=288690 $Y=211920
X878 1 2 4 ICV_13 $T=293940 187680 0 0 $X=293750 $Y=187440
X879 1 2 247 ICV_13 $T=300840 193120 0 0 $X=300650 $Y=192880
X880 1 2 256 ICV_13 $T=310500 198560 0 0 $X=310310 $Y=198320
X881 1 2 529 ICV_13 $T=311880 204000 1 0 $X=311690 $Y=201040
X882 1 2 258 ICV_13 $T=314640 209440 0 0 $X=314450 $Y=209200
X883 1 2 4 ICV_13 $T=322920 214880 0 0 $X=322730 $Y=214640
X884 1 2 536 ICV_13 $T=324760 214880 1 0 $X=324570 $Y=211920
X885 1 2 261 ICV_13 $T=327060 198560 0 0 $X=326870 $Y=198320
X886 1 2 ICV_14 $T=19780 176800 1 0 $X=19590 $Y=173840
X887 1 2 ICV_14 $T=33580 182240 0 0 $X=33390 $Y=182000
X888 1 2 ICV_14 $T=33580 198560 0 0 $X=33390 $Y=198320
X889 1 2 ICV_14 $T=47840 193120 1 0 $X=47650 $Y=190160
X890 1 2 ICV_14 $T=61640 209440 0 0 $X=61450 $Y=209200
X891 1 2 ICV_14 $T=75900 187680 1 0 $X=75710 $Y=184720
X892 1 2 ICV_14 $T=89700 204000 0 0 $X=89510 $Y=203760
X893 1 2 ICV_14 $T=117760 176800 0 0 $X=117570 $Y=176560
X894 1 2 ICV_14 $T=117760 204000 0 0 $X=117570 $Y=203760
X895 1 2 ICV_14 $T=117760 214880 0 0 $X=117570 $Y=214640
X896 1 2 ICV_14 $T=132020 193120 1 0 $X=131830 $Y=190160
X897 1 2 ICV_14 $T=132020 204000 1 0 $X=131830 $Y=201040
X898 1 2 ICV_14 $T=132020 209440 1 0 $X=131830 $Y=206480
X899 1 2 ICV_14 $T=145820 187680 0 0 $X=145630 $Y=187440
X900 1 2 ICV_14 $T=145820 204000 0 0 $X=145630 $Y=203760
X901 1 2 ICV_14 $T=201940 182240 0 0 $X=201750 $Y=182000
X902 1 2 ICV_14 $T=216200 182240 1 0 $X=216010 $Y=179280
X903 1 2 ICV_14 $T=244260 204000 1 0 $X=244070 $Y=201040
X904 1 2 ICV_14 $T=272320 182240 1 0 $X=272130 $Y=179280
X905 1 2 ICV_14 $T=286120 187680 0 0 $X=285930 $Y=187440
X906 1 2 ICV_14 $T=286120 204000 0 0 $X=285930 $Y=203760
X907 1 2 ICV_14 $T=314180 214880 0 0 $X=313990 $Y=214640
X908 1 14 ICV_15 $T=31740 176800 0 0 $X=31550 $Y=176560
X909 1 390 ICV_15 $T=31740 209440 0 0 $X=31550 $Y=209200
X910 1 28 ICV_15 $T=46000 198560 1 0 $X=45810 $Y=195600
X911 1 394 ICV_15 $T=46000 204000 1 0 $X=45810 $Y=201040
X912 1 50 ICV_15 $T=59800 176800 0 0 $X=59610 $Y=176560
X913 1 51 ICV_15 $T=59800 214880 0 0 $X=59610 $Y=214640
X914 1 65 ICV_15 $T=87860 193120 0 0 $X=87670 $Y=192880
X915 1 396 ICV_15 $T=87860 198560 0 0 $X=87670 $Y=198320
X916 1 396 ICV_15 $T=87860 209440 0 0 $X=87670 $Y=209200
X917 1 424 ICV_15 $T=102120 198560 1 0 $X=101930 $Y=195600
X918 1 426 ICV_15 $T=102120 204000 1 0 $X=101930 $Y=201040
X919 1 4 ICV_15 $T=115920 182240 0 0 $X=115730 $Y=182000
X920 1 429 ICV_15 $T=115920 193120 0 0 $X=115730 $Y=192880
X921 1 94 ICV_15 $T=130180 214880 1 0 $X=129990 $Y=211920
X922 1 4 ICV_15 $T=143980 182240 0 0 $X=143790 $Y=182000
X923 1 119 ICV_15 $T=143980 214880 0 0 $X=143790 $Y=214640
X924 1 461 ICV_15 $T=172040 176800 0 0 $X=171850 $Y=176560
X925 1 133 ICV_15 $T=172040 198560 0 0 $X=171850 $Y=198320
X926 1 170 ICV_15 $T=200100 187680 0 0 $X=199910 $Y=187440
X927 1 171 ICV_15 $T=200100 198560 0 0 $X=199910 $Y=198320
X928 1 475 ICV_15 $T=214360 209440 1 0 $X=214170 $Y=206480
X929 1 183 ICV_15 $T=214360 214880 1 0 $X=214170 $Y=211920
X930 1 4 ICV_15 $T=228160 193120 0 0 $X=227970 $Y=192880
X931 1 186 ICV_15 $T=228160 209440 0 0 $X=227970 $Y=209200
X932 1 490 ICV_15 $T=242420 209440 1 0 $X=242230 $Y=206480
X933 1 491 ICV_15 $T=242420 214880 1 0 $X=242230 $Y=211920
X934 1 212 ICV_15 $T=256220 176800 0 0 $X=256030 $Y=176560
X935 1 4 ICV_15 $T=256220 193120 0 0 $X=256030 $Y=192880
X936 1 220 ICV_15 $T=270480 187680 1 0 $X=270290 $Y=184720
X937 1 503 ICV_15 $T=270480 193120 1 0 $X=270290 $Y=190160
X938 1 172 ICV_15 $T=270480 214880 1 0 $X=270290 $Y=211920
X939 1 519 ICV_15 $T=298540 193120 1 0 $X=298350 $Y=190160
X940 1 4 ICV_15 $T=312340 187680 0 0 $X=312150 $Y=187440
X941 1 528 ICV_15 $T=312340 204000 0 0 $X=312150 $Y=203760
X942 1 2 374 ICV_16 $T=10120 182240 1 0 $X=9930 $Y=179280
X943 1 2 371 ICV_16 $T=11500 187680 1 0 $X=11310 $Y=184720
X944 1 2 372 ICV_16 $T=11500 193120 1 0 $X=11310 $Y=190160
X945 1 2 381 ICV_16 $T=24840 209440 1 0 $X=24650 $Y=206480
X946 1 2 32 ICV_16 $T=41400 187680 1 0 $X=41210 $Y=184720
X947 1 2 74 ICV_16 $T=81880 214880 0 0 $X=81690 $Y=214640
X948 1 2 72 ICV_16 $T=82800 176800 0 0 $X=82610 $Y=176560
X949 1 2 421 ICV_16 $T=95220 214880 1 0 $X=95030 $Y=211920
X950 1 2 85 ICV_16 $T=105340 204000 0 0 $X=105150 $Y=203760
X951 1 2 88 ICV_16 $T=109940 209440 0 0 $X=109750 $Y=209200
X952 1 2 98 ICV_16 $T=123740 193120 1 0 $X=123550 $Y=190160
X953 1 2 441 ICV_16 $T=137080 204000 1 0 $X=136890 $Y=201040
X954 1 2 447 ICV_16 $T=148580 193120 1 0 $X=148390 $Y=190160
X955 1 2 124 ICV_16 $T=150880 182240 1 0 $X=150690 $Y=179280
X956 1 2 126 ICV_16 $T=152260 198560 0 0 $X=152070 $Y=198320
X957 1 2 444 ICV_16 $T=153180 214880 1 0 $X=152990 $Y=211920
X958 1 2 446 ICV_16 $T=159620 204000 0 0 $X=159430 $Y=203760
X959 1 2 450 ICV_16 $T=161460 182240 1 0 $X=161270 $Y=179280
X960 1 2 129 ICV_16 $T=161920 176800 1 0 $X=161730 $Y=173840
X961 1 2 458 ICV_16 $T=181700 193120 1 0 $X=181510 $Y=190160
X962 1 2 144 ICV_16 $T=183080 204000 0 0 $X=182890 $Y=203760
X963 1 2 83 ICV_16 $T=185380 198560 0 0 $X=185190 $Y=198320
X964 1 2 76 ICV_16 $T=188600 193120 0 0 $X=188410 $Y=192880
X965 1 2 467 ICV_16 $T=189520 182240 1 0 $X=189330 $Y=179280
X966 1 2 151 ICV_16 $T=191820 204000 0 0 $X=191630 $Y=203760
X967 1 2 172 ICV_16 $T=203320 204000 0 0 $X=203130 $Y=203760
X968 1 2 215 ICV_16 $T=260820 176800 1 0 $X=260630 $Y=173840
X969 1 2 223 ICV_16 $T=273700 209440 1 0 $X=273510 $Y=206480
X970 1 2 228 ICV_16 $T=278760 204000 1 0 $X=278570 $Y=201040
X971 1 2 503 ICV_16 $T=280140 182240 1 0 $X=279950 $Y=179280
X972 1 2 245 ICV_16 $T=302220 204000 0 0 $X=302030 $Y=203760
X973 1 2 15 2 18 1 sky130_fd_sc_hd__inv_8 $T=21160 182240 1 0 $X=20970 $Y=179280
X974 1 2 373 2 380 1 sky130_fd_sc_hd__inv_8 $T=21160 198560 0 0 $X=20970 $Y=198320
X975 1 2 370 2 382 1 sky130_fd_sc_hd__inv_8 $T=23460 214880 0 0 $X=23270 $Y=214640
X976 1 2 32 2 395 1 sky130_fd_sc_hd__inv_8 $T=38640 187680 0 0 $X=38450 $Y=187440
X977 1 2 36 2 394 1 sky130_fd_sc_hd__inv_8 $T=41860 204000 0 0 $X=41670 $Y=203760
X978 1 2 38 2 388 1 sky130_fd_sc_hd__inv_8 $T=43240 176800 0 0 $X=43050 $Y=176560
X979 1 2 56 2 400 1 sky130_fd_sc_hd__inv_8 $T=63020 187680 0 0 $X=62830 $Y=187440
X980 1 2 58 2 407 1 sky130_fd_sc_hd__inv_8 $T=67620 198560 0 0 $X=67430 $Y=198320
X981 1 2 70 2 405 1 sky130_fd_sc_hd__inv_8 $T=77280 214880 1 0 $X=77090 $Y=211920
X982 1 2 72 2 75 1 sky130_fd_sc_hd__inv_8 $T=82800 182240 1 0 $X=82610 $Y=179280
X983 1 2 79 2 413 1 sky130_fd_sc_hd__inv_8 $T=92920 187680 1 0 $X=92730 $Y=184720
X984 1 2 426 2 419 1 sky130_fd_sc_hd__inv_8 $T=105340 204000 1 0 $X=105150 $Y=201040
X985 1 2 85 2 414 1 sky130_fd_sc_hd__inv_8 $T=105340 209440 1 0 $X=105150 $Y=206480
X986 1 2 88 2 425 1 sky130_fd_sc_hd__inv_8 $T=105340 214880 1 0 $X=105150 $Y=211920
X987 1 2 89 2 91 1 sky130_fd_sc_hd__inv_8 $T=109480 176800 0 0 $X=109290 $Y=176560
X988 1 2 98 2 436 1 sky130_fd_sc_hd__inv_8 $T=123740 193120 0 0 $X=123550 $Y=192880
X989 1 2 371 2 433 1 sky130_fd_sc_hd__inv_8 $T=127420 198560 0 0 $X=127230 $Y=198320
X990 1 2 103 2 112 1 sky130_fd_sc_hd__inv_8 $T=132480 182240 0 0 $X=132290 $Y=182000
X991 1 2 117 2 114 1 sky130_fd_sc_hd__inv_8 $T=141680 187680 1 0 $X=141490 $Y=184720
X992 1 2 126 2 443 1 sky130_fd_sc_hd__inv_8 $T=152260 204000 1 0 $X=152070 $Y=201040
X993 1 2 127 2 128 1 sky130_fd_sc_hd__inv_8 $T=155480 176800 0 0 $X=155290 $Y=176560
X994 1 2 449 2 123 1 sky130_fd_sc_hd__inv_8 $T=160540 182240 0 0 $X=160350 $Y=182000
X995 1 2 131 2 459 1 sky130_fd_sc_hd__inv_8 $T=168360 182240 1 0 $X=168170 $Y=179280
X996 1 2 133 2 458 1 sky130_fd_sc_hd__inv_8 $T=174800 204000 1 0 $X=174610 $Y=201040
X997 1 2 136 2 466 1 sky130_fd_sc_hd__inv_8 $T=175260 204000 0 0 $X=175070 $Y=203760
X998 1 2 145 2 465 1 sky130_fd_sc_hd__inv_8 $T=180320 176800 1 0 $X=180130 $Y=173840
X999 1 2 169 2 149 1 sky130_fd_sc_hd__inv_8 $T=197800 176800 1 0 $X=197610 $Y=173840
X1000 1 2 167 2 173 1 sky130_fd_sc_hd__inv_8 $T=203320 214880 0 0 $X=203130 $Y=214640
X1001 1 2 170 2 472 1 sky130_fd_sc_hd__inv_8 $T=204700 193120 1 0 $X=204510 $Y=190160
X1002 1 2 179 2 474 1 sky130_fd_sc_hd__inv_8 $T=212520 204000 0 0 $X=212330 $Y=203760
X1003 1 2 188 2 187 1 sky130_fd_sc_hd__inv_8 $T=217580 176800 1 0 $X=217390 $Y=173840
X1004 1 2 190 2 191 1 sky130_fd_sc_hd__inv_8 $T=222180 182240 0 0 $X=221990 $Y=182000
X1005 1 2 198 2 480 1 sky130_fd_sc_hd__inv_8 $T=234600 193120 1 0 $X=234410 $Y=190160
X1006 1 2 199 2 484 1 sky130_fd_sc_hd__inv_8 $T=235060 204000 1 0 $X=234870 $Y=201040
X1007 1 2 205 2 490 1 sky130_fd_sc_hd__inv_8 $T=246560 204000 1 0 $X=246370 $Y=201040
X1008 1 2 495 2 200 1 sky130_fd_sc_hd__inv_8 $T=248860 182240 0 0 $X=248670 $Y=182000
X1009 1 2 216 2 493 1 sky130_fd_sc_hd__inv_8 $T=258980 198560 1 0 $X=258790 $Y=195600
X1010 1 2 212 2 201 1 sky130_fd_sc_hd__inv_8 $T=259440 176800 0 0 $X=259250 $Y=176560
X1011 1 2 217 2 213 1 sky130_fd_sc_hd__inv_8 $T=264960 204000 0 0 $X=264770 $Y=203760
X1012 1 2 223 2 227 1 sky130_fd_sc_hd__inv_8 $T=273700 214880 1 0 $X=273510 $Y=211920
X1013 1 2 225 2 503 1 sky130_fd_sc_hd__inv_8 $T=275080 182240 1 0 $X=274890 $Y=179280
X1014 1 2 228 2 505 1 sky130_fd_sc_hd__inv_8 $T=277380 198560 0 0 $X=277190 $Y=198320
X1015 1 2 240 2 241 1 sky130_fd_sc_hd__inv_8 $T=292560 209440 1 0 $X=292370 $Y=206480
X1016 1 2 242 2 229 1 sky130_fd_sc_hd__inv_8 $T=301760 209440 0 0 $X=301570 $Y=209200
X1017 1 2 247 2 515 1 sky130_fd_sc_hd__inv_8 $T=304520 193120 0 0 $X=304330 $Y=192880
X1018 1 2 257 2 520 1 sky130_fd_sc_hd__inv_8 $T=314640 182240 1 0 $X=314450 $Y=179280
X1019 1 2 530 2 517 1 sky130_fd_sc_hd__inv_8 $T=315100 193120 1 0 $X=314910 $Y=190160
X1020 1 2 372 2 528 1 sky130_fd_sc_hd__inv_8 $T=315560 193120 0 0 $X=315370 $Y=192880
X1021 1 2 261 2 533 1 sky130_fd_sc_hd__inv_8 $T=330740 198560 0 0 $X=330550 $Y=198320
X1022 1 2 13 378 2 374 1 sky130_fd_sc_hd__nor2_4 $T=21160 176800 0 0 $X=20970 $Y=176560
X1023 1 2 14 375 2 376 1 sky130_fd_sc_hd__nor2_4 $T=21160 187680 0 0 $X=20970 $Y=187440
X1024 1 2 16 381 2 377 1 sky130_fd_sc_hd__nor2_4 $T=23000 209440 0 0 $X=22810 $Y=209200
X1025 1 2 16 383 2 384 1 sky130_fd_sc_hd__nor2_4 $T=28980 187680 1 0 $X=28790 $Y=184720
X1026 1 2 14 385 2 393 1 sky130_fd_sc_hd__nor2_4 $T=31740 204000 1 0 $X=31550 $Y=201040
X1027 1 2 14 391 2 31 1 sky130_fd_sc_hd__nor2_4 $T=34960 176800 0 0 $X=34770 $Y=176560
X1028 1 2 396 398 2 41 1 sky130_fd_sc_hd__nor2_4 $T=46920 214880 0 0 $X=46730 $Y=214640
X1029 1 2 396 399 2 402 1 sky130_fd_sc_hd__nor2_4 $T=53820 193120 0 0 $X=53630 $Y=192880
X1030 1 2 396 406 2 403 1 sky130_fd_sc_hd__nor2_4 $T=64400 198560 1 0 $X=64210 $Y=195600
X1031 1 2 60 63 2 408 1 sky130_fd_sc_hd__nor2_4 $T=68080 176800 1 0 $X=67890 $Y=173840
X1032 1 2 73 411 2 410 1 sky130_fd_sc_hd__nor2_4 $T=81420 198560 1 0 $X=81230 $Y=195600
X1033 1 2 396 417 2 420 1 sky130_fd_sc_hd__nor2_4 $T=91080 198560 0 0 $X=90890 $Y=198320
X1034 1 2 396 418 2 421 1 sky130_fd_sc_hd__nor2_4 $T=91080 209440 0 0 $X=90890 $Y=209200
X1035 1 2 73 415 2 423 1 sky130_fd_sc_hd__nor2_4 $T=92460 209440 1 0 $X=92270 $Y=206480
X1036 1 2 90 428 2 427 1 sky130_fd_sc_hd__nor2_4 $T=114080 209440 1 0 $X=113890 $Y=206480
X1037 1 2 90 432 2 429 1 sky130_fd_sc_hd__nor2_4 $T=119600 198560 0 0 $X=119410 $Y=198320
X1038 1 2 99 431 2 430 1 sky130_fd_sc_hd__nor2_4 $T=123740 176800 0 0 $X=123550 $Y=176560
X1039 1 2 99 438 2 440 1 sky130_fd_sc_hd__nor2_4 $T=133400 182240 1 0 $X=133210 $Y=179280
X1040 1 2 439 111 2 441 1 sky130_fd_sc_hd__nor2_4 $T=136160 214880 1 0 $X=135970 $Y=211920
X1041 1 2 102 442 2 447 1 sky130_fd_sc_hd__nor2_4 $T=145820 182240 1 0 $X=145630 $Y=179280
X1042 1 2 102 124 2 445 1 sky130_fd_sc_hd__nor2_4 $T=147660 176800 0 0 $X=147470 $Y=176560
X1043 1 2 90 446 2 448 1 sky130_fd_sc_hd__nor2_4 $T=151340 209440 1 0 $X=151150 $Y=206480
X1044 1 2 130 453 2 450 1 sky130_fd_sc_hd__nor2_4 $T=166060 187680 0 0 $X=165870 $Y=187440
X1045 1 2 130 454 2 451 1 sky130_fd_sc_hd__nor2_4 $T=166060 193120 0 0 $X=165870 $Y=192880
X1046 1 2 137 457 2 452 1 sky130_fd_sc_hd__nor2_4 $T=172500 209440 1 0 $X=172310 $Y=206480
X1047 1 2 130 463 2 141 1 sky130_fd_sc_hd__nor2_4 $T=177560 176800 0 0 $X=177370 $Y=176560
X1048 1 2 174 470 2 468 1 sky130_fd_sc_hd__nor2_4 $T=207000 187680 0 0 $X=206810 $Y=187440
X1049 1 2 178 473 2 471 1 sky130_fd_sc_hd__nor2_4 $T=208380 204000 1 0 $X=208190 $Y=201040
X1050 1 2 174 479 2 476 1 sky130_fd_sc_hd__nor2_4 $T=218500 182240 1 0 $X=218310 $Y=179280
X1051 1 2 178 477 2 481 1 sky130_fd_sc_hd__nor2_4 $T=222180 198560 0 0 $X=221990 $Y=198320
X1052 1 2 178 482 2 483 1 sky130_fd_sc_hd__nor2_4 $T=231380 198560 0 0 $X=231190 $Y=198320
X1053 1 2 174 487 2 492 1 sky130_fd_sc_hd__nor2_4 $T=240120 182240 0 0 $X=239930 $Y=182000
X1054 1 2 202 488 2 489 1 sky130_fd_sc_hd__nor2_4 $T=242880 204000 0 0 $X=242690 $Y=203760
X1055 1 2 204 206 2 497 1 sky130_fd_sc_hd__nor2_4 $T=247480 176800 0 0 $X=247290 $Y=176560
X1056 1 2 202 496 2 498 1 sky130_fd_sc_hd__nor2_4 $T=250700 198560 1 0 $X=250510 $Y=195600
X1057 1 2 202 499 2 500 1 sky130_fd_sc_hd__nor2_4 $T=258980 209440 1 0 $X=258790 $Y=206480
X1058 1 2 439 501 2 502 1 sky130_fd_sc_hd__nor2_4 $T=269100 187680 0 0 $X=268910 $Y=187440
X1059 1 2 439 506 2 504 1 sky130_fd_sc_hd__nor2_4 $T=273700 204000 1 0 $X=273510 $Y=201040
X1060 1 2 222 232 2 511 1 sky130_fd_sc_hd__nor2_4 $T=284740 214880 1 0 $X=284550 $Y=211920
X1061 1 2 230 514 2 518 1 sky130_fd_sc_hd__nor2_4 $T=289340 182240 0 0 $X=289150 $Y=182000
X1062 1 2 222 236 2 516 1 sky130_fd_sc_hd__nor2_4 $T=292560 214880 1 0 $X=292370 $Y=211920
X1063 1 2 439 522 2 524 1 sky130_fd_sc_hd__nor2_4 $T=301760 187680 1 0 $X=301570 $Y=184720
X1064 1 2 439 519 2 525 1 sky130_fd_sc_hd__nor2_4 $T=301760 193120 1 0 $X=301570 $Y=190160
X1065 1 2 252 526 2 527 1 sky130_fd_sc_hd__nor2_4 $T=307740 204000 1 0 $X=307550 $Y=201040
X1066 1 2 252 534 2 535 1 sky130_fd_sc_hd__nor2_4 $T=320620 209440 0 0 $X=320430 $Y=209200
X1067 1 2 252 531 2 536 1 sky130_fd_sc_hd__nor2_4 $T=320620 214880 1 0 $X=320430 $Y=211920
X1068 1 2 18 19 22 21 2 378 1 sky130_fd_sc_hd__o22a_4 $T=22540 176800 1 0 $X=22350 $Y=173840
X1069 1 2 380 20 17 379 2 375 1 sky130_fd_sc_hd__o22a_4 $T=23460 193120 0 0 $X=23270 $Y=192880
X1070 1 2 382 23 390 386 2 381 1 sky130_fd_sc_hd__o22a_4 $T=34500 214880 1 0 $X=34310 $Y=211920
X1071 1 2 27 23 390 35 2 29 1 sky130_fd_sc_hd__o22a_4 $T=34960 214880 0 0 $X=34770 $Y=214640
X1072 1 2 388 20 17 392 2 391 1 sky130_fd_sc_hd__o22a_4 $T=35880 182240 0 0 $X=35690 $Y=182000
X1073 1 2 395 23 390 389 2 383 1 sky130_fd_sc_hd__o22a_4 $T=35880 198560 1 0 $X=35690 $Y=195600
X1074 1 2 394 20 17 387 2 385 1 sky130_fd_sc_hd__o22a_4 $T=35880 198560 0 0 $X=35690 $Y=198320
X1075 1 2 44 23 390 397 2 398 1 sky130_fd_sc_hd__o22a_4 $T=49220 214880 1 0 $X=49030 $Y=211920
X1076 1 2 400 23 390 401 2 399 1 sky130_fd_sc_hd__o22a_4 $T=54280 198560 1 0 $X=54090 $Y=195600
X1077 1 2 405 51 66 59 2 53 1 sky130_fd_sc_hd__o22a_4 $T=68080 214880 0 0 $X=67890 $Y=214640
X1078 1 2 407 65 64 409 2 406 1 sky130_fd_sc_hd__o22a_4 $T=73140 193120 0 0 $X=72950 $Y=192880
X1079 1 2 75 65 64 77 2 63 1 sky130_fd_sc_hd__o22a_4 $T=79120 176800 1 0 $X=78930 $Y=173840
X1080 1 2 413 80 78 416 2 411 1 sky130_fd_sc_hd__o22a_4 $T=90160 193120 1 0 $X=89970 $Y=190160
X1081 1 2 414 65 64 412 2 418 1 sky130_fd_sc_hd__o22a_4 $T=90160 204000 1 0 $X=89970 $Y=201040
X1082 1 2 419 65 64 422 2 417 1 sky130_fd_sc_hd__o22a_4 $T=91080 198560 1 0 $X=90890 $Y=195600
X1083 1 2 425 80 78 424 2 415 1 sky130_fd_sc_hd__o22a_4 $T=96600 193120 0 0 $X=96410 $Y=192880
X1084 1 2 433 95 94 434 2 428 1 sky130_fd_sc_hd__o22a_4 $T=121900 209440 1 0 $X=121710 $Y=206480
X1085 1 2 436 95 94 435 2 432 1 sky130_fd_sc_hd__o22a_4 $T=124200 204000 0 0 $X=124010 $Y=203760
X1086 1 2 112 113 109 115 2 431 1 sky130_fd_sc_hd__o22a_4 $T=133400 176800 1 0 $X=133210 $Y=173840
X1087 1 2 110 95 437 94 2 108 1 sky130_fd_sc_hd__o22a_4 $T=133860 214880 0 0 $X=133670 $Y=214640
X1088 1 2 114 113 109 105 2 438 1 sky130_fd_sc_hd__o22a_4 $T=135700 176800 0 0 $X=135510 $Y=176560
X1089 1 2 123 113 109 125 2 442 1 sky130_fd_sc_hd__o22a_4 $T=146740 176800 1 0 $X=146550 $Y=173840
X1090 1 2 443 95 94 444 2 446 1 sky130_fd_sc_hd__o22a_4 $T=147200 209440 0 0 $X=147010 $Y=209200
X1091 1 2 459 460 462 456 2 453 1 sky130_fd_sc_hd__o22a_4 $T=174800 187680 1 0 $X=174610 $Y=184720
X1092 1 2 458 460 462 455 2 454 1 sky130_fd_sc_hd__o22a_4 $T=175260 193120 0 0 $X=175070 $Y=192880
X1093 1 2 466 460 462 464 2 457 1 sky130_fd_sc_hd__o22a_4 $T=176180 198560 1 0 $X=175990 $Y=195600
X1094 1 2 465 460 462 461 2 463 1 sky130_fd_sc_hd__o22a_4 $T=178020 182240 1 0 $X=177830 $Y=179280
X1095 1 2 149 460 462 467 2 150 1 sky130_fd_sc_hd__o22a_4 $T=186300 176800 0 0 $X=186110 $Y=176560
X1096 1 2 472 50 52 469 2 470 1 sky130_fd_sc_hd__o22a_4 $T=205620 187680 1 0 $X=205430 $Y=184720
X1097 1 2 177 183 182 185 2 180 1 sky130_fd_sc_hd__o22a_4 $T=210680 214880 0 0 $X=210490 $Y=214640
X1098 1 2 474 183 182 475 2 473 1 sky130_fd_sc_hd__o22a_4 $T=217580 209440 1 0 $X=217390 $Y=206480
X1099 1 2 480 183 182 478 2 482 1 sky130_fd_sc_hd__o22a_4 $T=223560 204000 1 0 $X=223370 $Y=201040
X1100 1 2 191 196 197 193 2 479 1 sky130_fd_sc_hd__o22a_4 $T=225860 176800 1 0 $X=225670 $Y=173840
X1101 1 2 484 183 182 485 2 477 1 sky130_fd_sc_hd__o22a_4 $T=226780 209440 1 0 $X=226590 $Y=206480
X1102 1 2 200 196 197 486 2 487 1 sky130_fd_sc_hd__o22a_4 $T=237360 176800 0 0 $X=237170 $Y=176560
X1103 1 2 490 207 203 491 2 488 1 sky130_fd_sc_hd__o22a_4 $T=247020 209440 0 0 $X=246830 $Y=209200
X1104 1 2 493 207 203 494 2 496 1 sky130_fd_sc_hd__o22a_4 $T=248860 209440 1 0 $X=248670 $Y=206480
X1105 1 2 213 207 203 214 2 499 1 sky130_fd_sc_hd__o22a_4 $T=254840 214880 1 0 $X=254650 $Y=211920
X1106 1 2 503 509 510 507 2 501 1 sky130_fd_sc_hd__o22a_4 $T=278760 187680 1 0 $X=278570 $Y=184720
X1107 1 2 505 509 510 508 2 506 1 sky130_fd_sc_hd__o22a_4 $T=280140 193120 1 0 $X=279950 $Y=190160
X1108 1 2 515 509 510 513 2 514 1 sky130_fd_sc_hd__o22a_4 $T=290260 187680 1 0 $X=290070 $Y=184720
X1109 1 2 517 509 510 512 2 519 1 sky130_fd_sc_hd__o22a_4 $T=294400 193120 0 0 $X=294210 $Y=192880
X1110 1 2 520 509 510 521 2 522 1 sky130_fd_sc_hd__o22a_4 $T=298080 182240 0 0 $X=297890 $Y=182000
X1111 1 2 249 246 248 523 2 255 1 sky130_fd_sc_hd__o22a_4 $T=310500 214880 1 0 $X=310310 $Y=211920
X1112 1 2 528 246 248 529 2 526 1 sky130_fd_sc_hd__o22a_4 $T=313720 209440 1 0 $X=313530 $Y=206480
X1113 1 2 258 246 248 259 2 531 1 sky130_fd_sc_hd__o22a_4 $T=316480 214880 0 0 $X=316290 $Y=214640
X1114 1 2 533 246 248 532 2 534 1 sky130_fd_sc_hd__o22a_4 $T=321540 204000 0 0 $X=321350 $Y=203760
X1115 1 2 33 2 14 1 sky130_fd_sc_hd__buf_1 $T=39100 187680 1 0 $X=38910 $Y=184720
X1116 1 2 33 2 16 1 sky130_fd_sc_hd__buf_1 $T=41400 193120 1 0 $X=41210 $Y=190160
X1117 1 2 40 2 20 1 sky130_fd_sc_hd__buf_1 $T=46460 182240 0 0 $X=46270 $Y=182000
X1118 1 2 42 2 17 1 sky130_fd_sc_hd__buf_1 $T=49220 187680 1 0 $X=49030 $Y=184720
X1119 1 2 43 2 24 1 sky130_fd_sc_hd__buf_1 $T=49680 187680 0 0 $X=49490 $Y=187440
X1120 1 2 40 2 23 1 sky130_fd_sc_hd__buf_1 $T=50600 193120 1 0 $X=50410 $Y=190160
X1121 1 2 43 2 28 1 sky130_fd_sc_hd__buf_1 $T=51060 176800 1 0 $X=50870 $Y=173840
X1122 1 2 42 2 390 1 sky130_fd_sc_hd__buf_1 $T=54740 187680 0 0 $X=54550 $Y=187440
X1123 1 2 39 2 48 1 sky130_fd_sc_hd__buf_1 $T=56580 209440 0 0 $X=56390 $Y=209200
X1124 1 2 34 2 49 1 sky130_fd_sc_hd__buf_1 $T=57040 193120 1 0 $X=56850 $Y=190160
X1125 1 2 52 2 22 1 sky130_fd_sc_hd__buf_1 $T=62100 182240 1 0 $X=61910 $Y=179280
X1126 1 2 33 2 396 1 sky130_fd_sc_hd__buf_1 $T=62100 193120 1 0 $X=61910 $Y=190160
X1127 1 2 50 2 19 1 sky130_fd_sc_hd__buf_1 $T=63020 176800 0 0 $X=62830 $Y=176560
X1128 1 2 26 2 54 1 sky130_fd_sc_hd__buf_1 $T=63020 214880 0 0 $X=62830 $Y=214640
X1129 1 2 50 2 51 1 sky130_fd_sc_hd__buf_1 $T=74060 204000 0 0 $X=73870 $Y=203760
X1130 1 2 52 2 66 1 sky130_fd_sc_hd__buf_1 $T=75900 198560 0 0 $X=75710 $Y=198320
X1131 1 2 67 2 57 1 sky130_fd_sc_hd__buf_1 $T=77280 209440 1 0 $X=77090 $Y=206480
X1132 1 2 67 2 73 1 sky130_fd_sc_hd__buf_1 $T=80500 204000 1 0 $X=80310 $Y=201040
X1133 1 2 76 2 62 1 sky130_fd_sc_hd__buf_1 $T=83260 209440 0 0 $X=83070 $Y=209200
X1134 1 2 40 2 65 1 sky130_fd_sc_hd__buf_1 $T=83720 182240 0 0 $X=83530 $Y=182000
X1135 1 2 42 2 64 1 sky130_fd_sc_hd__buf_1 $T=90620 182240 1 0 $X=90430 $Y=179280
X1136 1 2 76 2 82 1 sky130_fd_sc_hd__buf_1 $T=92000 204000 0 0 $X=91810 $Y=203760
X1137 1 2 50 2 80 1 sky130_fd_sc_hd__buf_1 $T=96600 176800 0 0 $X=96410 $Y=176560
X1138 1 2 52 2 78 1 sky130_fd_sc_hd__buf_1 $T=98440 182240 0 0 $X=98250 $Y=182000
X1139 1 2 84 2 404 1 sky130_fd_sc_hd__buf_1 $T=98900 182240 1 0 $X=98710 $Y=179280
X1140 1 2 92 2 93 1 sky130_fd_sc_hd__buf_1 $T=119600 209440 0 0 $X=119410 $Y=209200
X1141 1 2 33 2 99 1 sky130_fd_sc_hd__buf_1 $T=124200 182240 1 0 $X=124010 $Y=179280
X1142 1 2 67 2 102 1 sky130_fd_sc_hd__buf_1 $T=126960 176800 1 0 $X=126770 $Y=173840
X1143 1 2 104 2 106 1 sky130_fd_sc_hd__buf_1 $T=129260 187680 0 0 $X=129070 $Y=187440
X1144 1 2 120 2 439 1 sky130_fd_sc_hd__buf_1 $T=145360 198560 1 0 $X=145170 $Y=195600
X1145 1 2 122 2 94 1 sky130_fd_sc_hd__buf_1 $T=149960 214880 0 0 $X=149770 $Y=214640
X1146 1 2 52 2 134 1 sky130_fd_sc_hd__buf_1 $T=171120 176800 1 0 $X=170930 $Y=173840
X1147 1 2 83 2 146 1 sky130_fd_sc_hd__buf_1 $T=182620 204000 1 0 $X=182430 $Y=201040
X1148 1 2 144 2 137 1 sky130_fd_sc_hd__buf_1 $T=183080 209440 1 0 $X=182890 $Y=206480
X1149 1 2 144 2 148 1 sky130_fd_sc_hd__buf_1 $T=185380 209440 0 0 $X=185190 $Y=209200
X1150 1 2 151 2 462 1 sky130_fd_sc_hd__buf_1 $T=189520 193120 1 0 $X=189330 $Y=190160
X1151 1 2 76 2 116 1 sky130_fd_sc_hd__buf_1 $T=189520 198560 1 0 $X=189330 $Y=195600
X1152 1 2 153 2 460 1 sky130_fd_sc_hd__buf_1 $T=189980 187680 0 0 $X=189790 $Y=187440
X1153 1 2 151 2 155 1 sky130_fd_sc_hd__buf_1 $T=191820 209440 1 0 $X=191630 $Y=206480
X1154 1 2 81 2 156 1 sky130_fd_sc_hd__buf_1 $T=192280 198560 0 0 $X=192090 $Y=198320
X1155 1 2 69 2 162 1 sky130_fd_sc_hd__buf_1 $T=195040 193120 1 0 $X=194850 $Y=190160
X1156 1 2 159 2 120 1 sky130_fd_sc_hd__buf_1 $T=195040 198560 1 0 $X=194850 $Y=195600
X1157 1 2 163 2 164 1 sky130_fd_sc_hd__buf_1 $T=196420 176800 0 0 $X=196230 $Y=176560
X1158 1 2 158 2 165 1 sky130_fd_sc_hd__buf_1 $T=197340 182240 1 0 $X=197150 $Y=179280
X1159 1 2 171 2 90 1 sky130_fd_sc_hd__buf_1 $T=201020 204000 1 0 $X=200830 $Y=201040
X1160 1 2 166 2 118 1 sky130_fd_sc_hd__buf_1 $T=201940 198560 1 0 $X=201750 $Y=195600
X1161 1 2 172 2 97 1 sky130_fd_sc_hd__buf_1 $T=202400 209440 1 0 $X=202210 $Y=206480
X1162 1 2 176 2 159 1 sky130_fd_sc_hd__buf_1 $T=205620 176800 1 0 $X=205430 $Y=173840
X1163 1 2 171 2 178 1 sky130_fd_sc_hd__buf_1 $T=217580 204000 1 0 $X=217390 $Y=201040
X1164 1 2 122 2 182 1 sky130_fd_sc_hd__buf_1 $T=226780 214880 1 0 $X=226590 $Y=211920
X1165 1 2 172 2 186 1 sky130_fd_sc_hd__buf_1 $T=235060 214880 1 0 $X=234870 $Y=211920
X1166 1 2 122 2 203 1 sky130_fd_sc_hd__buf_1 $T=240580 214880 0 0 $X=240390 $Y=214640
X1167 1 2 171 2 202 1 sky130_fd_sc_hd__buf_1 $T=250700 204000 0 0 $X=250510 $Y=203760
X1168 1 2 172 2 210 1 sky130_fd_sc_hd__buf_1 $T=264960 214880 1 0 $X=264770 $Y=211920
X1169 1 2 172 2 221 1 sky130_fd_sc_hd__buf_1 $T=270480 214880 0 0 $X=270290 $Y=214640
X1170 1 2 120 2 224 1 sky130_fd_sc_hd__buf_1 $T=273700 187680 1 0 $X=273510 $Y=184720
X1171 1 2 120 2 230 1 sky130_fd_sc_hd__buf_1 $T=280140 176800 0 0 $X=279950 $Y=176560
X1172 1 2 120 2 233 1 sky130_fd_sc_hd__buf_1 $T=288880 176800 1 0 $X=288690 $Y=173840
X1173 1 2 237 2 220 1 sky130_fd_sc_hd__buf_1 $T=292100 176800 0 0 $X=291910 $Y=176560
X1174 1 2 238 2 509 1 sky130_fd_sc_hd__buf_1 $T=292100 193120 1 0 $X=291910 $Y=190160
X1175 1 2 239 2 510 1 sky130_fd_sc_hd__buf_1 $T=293940 182240 1 0 $X=293750 $Y=179280
X1176 1 2 244 2 246 1 sky130_fd_sc_hd__buf_1 $T=301760 214880 1 0 $X=301570 $Y=211920
X1177 1 2 245 2 248 1 sky130_fd_sc_hd__buf_1 $T=302220 209440 1 0 $X=302030 $Y=206480
X1178 1 2 25 380 28 2 379 1 sky130_fd_sc_hd__o21a_4 $T=34960 193120 0 0 $X=34770 $Y=192880
X1179 1 2 30 382 24 2 386 1 sky130_fd_sc_hd__o21a_4 $T=37260 209440 0 0 $X=37070 $Y=209200
X1180 1 2 34 388 28 2 392 1 sky130_fd_sc_hd__o21a_4 $T=38640 182240 1 0 $X=38450 $Y=179280
X1181 1 2 37 395 24 2 389 1 sky130_fd_sc_hd__o21a_4 $T=43240 193120 0 0 $X=43050 $Y=192880
X1182 1 2 39 394 28 2 387 1 sky130_fd_sc_hd__o21a_4 $T=46000 198560 0 0 $X=45810 $Y=198320
X1183 1 2 47 44 404 2 397 1 sky130_fd_sc_hd__o21a_4 $T=55200 209440 1 0 $X=55010 $Y=206480
X1184 1 2 55 400 404 2 401 1 sky130_fd_sc_hd__o21a_4 $T=63480 193120 0 0 $X=63290 $Y=192880
X1185 1 2 26 405 62 2 59 1 sky130_fd_sc_hd__o21a_4 $T=66700 214880 1 0 $X=66510 $Y=211920
X1186 1 2 69 407 404 2 409 1 sky130_fd_sc_hd__o21a_4 $T=77280 193120 1 0 $X=77090 $Y=190160
X1187 1 2 81 413 82 2 416 1 sky130_fd_sc_hd__o21a_4 $T=93840 187680 0 0 $X=93650 $Y=187440
X1188 1 2 83 425 82 2 424 1 sky130_fd_sc_hd__o21a_4 $T=98900 204000 0 0 $X=98710 $Y=203760
X1189 1 2 81 414 404 2 412 1 sky130_fd_sc_hd__o21a_4 $T=105340 198560 1 0 $X=105150 $Y=195600
X1190 1 2 83 419 404 2 422 1 sky130_fd_sc_hd__o21a_4 $T=106720 193120 0 0 $X=106530 $Y=192880
X1191 1 2 101 433 97 2 434 1 sky130_fd_sc_hd__o21a_4 $T=124660 209440 0 0 $X=124470 $Y=209200
X1192 1 2 106 436 97 2 435 1 sky130_fd_sc_hd__o21a_4 $T=134320 204000 0 0 $X=134130 $Y=203760
X1193 1 2 107 110 116 2 437 1 sky130_fd_sc_hd__o21a_4 $T=136620 209440 0 0 $X=136430 $Y=209200
X1194 1 2 118 443 97 2 444 1 sky130_fd_sc_hd__o21a_4 $T=146740 214880 1 0 $X=146550 $Y=211920
X1195 1 2 135 459 139 2 456 1 sky130_fd_sc_hd__o21a_4 $T=175260 187680 0 0 $X=175070 $Y=187440
X1196 1 2 142 458 139 2 455 1 sky130_fd_sc_hd__o21a_4 $T=175260 193120 1 0 $X=175070 $Y=190160
X1197 1 2 140 466 139 2 464 1 sky130_fd_sc_hd__o21a_4 $T=178940 198560 0 0 $X=178750 $Y=198320
X1198 1 2 143 465 139 2 461 1 sky130_fd_sc_hd__o21a_4 $T=182160 182240 0 0 $X=181970 $Y=182000
X1199 1 2 154 149 139 2 467 1 sky130_fd_sc_hd__o21a_4 $T=189520 176800 1 0 $X=189330 $Y=173840
X1200 1 2 175 472 116 2 469 1 sky130_fd_sc_hd__o21a_4 $T=206540 182240 0 0 $X=206350 $Y=182000
X1201 1 2 184 474 186 2 475 1 sky130_fd_sc_hd__o21a_4 $T=217580 214880 1 0 $X=217390 $Y=211920
X1202 1 2 49 480 186 2 478 1 sky130_fd_sc_hd__o21a_4 $T=220800 204000 0 0 $X=220610 $Y=203760
X1203 1 2 192 191 116 2 193 1 sky130_fd_sc_hd__o21a_4 $T=226320 182240 1 0 $X=226130 $Y=179280
X1204 1 2 194 484 186 2 485 1 sky130_fd_sc_hd__o21a_4 $T=231380 209440 0 0 $X=231190 $Y=209200
X1205 1 2 208 200 116 2 486 1 sky130_fd_sc_hd__o21a_4 $T=245640 176800 1 0 $X=245450 $Y=173840
X1206 1 2 54 493 186 2 494 1 sky130_fd_sc_hd__o21a_4 $T=245640 214880 1 0 $X=245450 $Y=211920
X1207 1 2 209 490 210 2 491 1 sky130_fd_sc_hd__o21a_4 $T=248860 214880 0 0 $X=248670 $Y=214640
X1208 1 2 162 503 220 2 507 1 sky130_fd_sc_hd__o21a_4 $T=276920 187680 0 0 $X=276730 $Y=187440
X1209 1 2 156 505 220 2 508 1 sky130_fd_sc_hd__o21a_4 $T=276920 193120 0 0 $X=276730 $Y=192880
X1210 1 2 146 229 210 2 226 1 sky130_fd_sc_hd__o21a_4 $T=276920 214880 0 0 $X=276730 $Y=214640
X1211 1 2 146 517 234 2 512 1 sky130_fd_sc_hd__o21a_4 $T=287960 204000 1 0 $X=287770 $Y=201040
X1212 1 2 165 515 220 2 513 1 sky130_fd_sc_hd__o21a_4 $T=288420 187680 0 0 $X=288230 $Y=187440
X1213 1 2 164 241 221 2 235 1 sky130_fd_sc_hd__o21a_4 $T=289800 214880 0 0 $X=289610 $Y=214640
X1214 1 2 164 520 220 2 521 1 sky130_fd_sc_hd__o21a_4 $T=301760 182240 1 0 $X=301570 $Y=179280
X1215 1 2 243 249 250 2 523 1 sky130_fd_sc_hd__o21a_4 $T=304980 214880 0 0 $X=304790 $Y=214640
X1216 1 2 256 528 250 2 529 1 sky130_fd_sc_hd__o21a_4 $T=315560 204000 1 0 $X=315370 $Y=201040
X1217 1 2 260 533 250 2 532 1 sky130_fd_sc_hd__o21a_4 $T=321540 198560 0 0 $X=321350 $Y=198320
X1218 1 2 4 ICV_22 $T=6900 182240 0 0 $X=6710 $Y=182000
X1219 1 2 379 ICV_22 $T=22080 187680 1 0 $X=21890 $Y=184720
X1220 1 2 30 ICV_22 $T=34040 209440 0 0 $X=33850 $Y=209200
X1221 1 2 46 ICV_22 $T=52440 176800 1 0 $X=52250 $Y=173840
X1222 1 2 67 ICV_22 $T=79120 198560 0 0 $X=78930 $Y=198320
X1223 1 2 4 ICV_22 $T=95220 198560 0 0 $X=95030 $Y=198320
X1224 1 2 4 ICV_22 $T=95220 209440 0 0 $X=95030 $Y=209200
X1225 1 2 92 ICV_22 $T=118220 209440 1 0 $X=118030 $Y=206480
X1226 1 2 117 ICV_22 $T=140300 182240 0 0 $X=140110 $Y=182000
X1227 1 2 102 ICV_22 $T=143520 176800 1 0 $X=143330 $Y=173840
X1228 1 2 90 ICV_22 $T=149040 204000 1 0 $X=148850 $Y=201040
X1229 1 2 130 ICV_22 $T=162840 187680 0 0 $X=162650 $Y=187440
X1230 1 2 130 ICV_22 $T=162840 193120 0 0 $X=162650 $Y=192880
X1231 1 2 462 ICV_22 $T=174340 176800 0 0 $X=174150 $Y=176560
X1232 1 2 210 ICV_22 $T=273700 214880 0 0 $X=273510 $Y=214640
X1233 1 2 165 ICV_22 $T=287040 187680 1 0 $X=286850 $Y=184720
X1234 1 2 252 ICV_22 $T=317400 209440 0 0 $X=317210 $Y=209200
X1235 1 2 250 ICV_22 $T=318320 198560 0 0 $X=318130 $Y=198320
X1236 1 2 248 ICV_22 $T=318320 204000 0 0 $X=318130 $Y=203760
X1237 1 2 535 ICV_22 $T=324760 193120 1 0 $X=324570 $Y=190160
X1238 1 2 ICV_23 $T=8740 204000 1 0 $X=8550 $Y=201040
X1239 1 2 ICV_23 $T=8740 204000 0 0 $X=8550 $Y=203760
X1240 1 2 ICV_23 $T=19780 204000 0 0 $X=19590 $Y=203760
X1241 1 2 ICV_23 $T=47380 176800 0 0 $X=47190 $Y=176560
X1242 1 2 ICV_23 $T=54740 176800 1 0 $X=54550 $Y=173840
X1243 1 2 ICV_23 $T=78660 209440 1 0 $X=78470 $Y=206480
X1244 1 2 ICV_23 $T=81420 214880 1 0 $X=81230 $Y=211920
X1245 1 2 ICV_23 $T=85560 176800 1 0 $X=85370 $Y=173840
X1246 1 2 ICV_23 $T=101200 187680 0 0 $X=101010 $Y=187440
X1247 1 2 ICV_23 $T=101660 182240 0 0 $X=101470 $Y=182000
X1248 1 2 ICV_23 $T=105800 214880 0 0 $X=105610 $Y=214640
X1249 1 2 ICV_23 $T=109940 193120 1 0 $X=109750 $Y=190160
X1250 1 2 ICV_23 $T=110400 176800 1 0 $X=110210 $Y=173840
X1251 1 2 ICV_23 $T=115460 187680 1 0 $X=115270 $Y=184720
X1252 1 2 ICV_23 $T=127880 193120 0 0 $X=127690 $Y=192880
X1253 1 2 ICV_23 $T=131560 198560 0 0 $X=131370 $Y=198320
X1254 1 2 ICV_23 $T=146740 198560 1 0 $X=146550 $Y=195600
X1255 1 2 ICV_23 $T=148120 193120 0 0 $X=147930 $Y=192880
X1256 1 2 ICV_23 $T=153180 214880 0 0 $X=152990 $Y=214640
X1257 1 2 ICV_23 $T=176640 214880 1 0 $X=176450 $Y=211920
X1258 1 2 ICV_23 $T=187680 182240 0 0 $X=187490 $Y=182000
X1259 1 2 ICV_23 $T=211140 187680 0 0 $X=210950 $Y=187440
X1260 1 2 ICV_23 $T=228160 187680 1 0 $X=227970 $Y=184720
X1261 1 2 ICV_23 $T=235520 187680 0 0 $X=235330 $Y=187440
X1262 1 2 ICV_23 $T=246560 187680 0 0 $X=246370 $Y=187440
X1263 1 2 ICV_23 $T=256220 187680 1 0 $X=256030 $Y=184720
X1264 1 2 ICV_23 $T=262200 198560 0 0 $X=262010 $Y=198320
X1265 1 2 ICV_23 $T=263580 176800 0 0 $X=263390 $Y=176560
X1266 1 2 ICV_23 $T=269100 204000 0 0 $X=268910 $Y=203760
X1267 1 2 ICV_23 $T=292560 198560 0 0 $X=292370 $Y=198320
X1268 1 2 ICV_23 $T=317400 187680 1 0 $X=317210 $Y=184720
X1269 1 2 ICV_23 $T=326600 209440 0 0 $X=326410 $Y=209200
X1270 1 2 ICV_23 $T=327980 204000 0 0 $X=327790 $Y=203760
X1271 1 2 ICV_23 $T=337640 214880 1 0 $X=337450 $Y=211920
X1272 1 2 391 31 ICV_27 $T=34040 176800 1 0 $X=33850 $Y=173840
X1273 1 2 392 17 ICV_27 $T=34040 182240 1 0 $X=33850 $Y=179280
X1274 1 2 4 393 ICV_27 $T=34960 204000 0 0 $X=34770 $Y=203760
X1275 1 2 24 382 ICV_27 $T=43700 209440 0 0 $X=43510 $Y=209200
X1276 1 2 4 403 ICV_27 $T=56580 198560 0 0 $X=56390 $Y=198320
X1277 1 2 34 42 ICV_27 $T=57040 187680 0 0 $X=56850 $Y=187440
X1278 1 2 4 410 ICV_27 $T=78660 182240 0 0 $X=78470 $Y=182000
X1279 1 2 4 87 ICV_27 $T=104420 176800 0 0 $X=104230 $Y=176560
X1280 1 2 4 432 ICV_27 $T=119140 193120 0 0 $X=118950 $Y=192880
X1281 1 2 94 94 ICV_27 $T=120060 214880 1 0 $X=119870 $Y=211920
X1282 1 2 462 460 ICV_27 $T=175260 182240 0 0 $X=175070 $Y=182000
X1283 1 2 157 161 ICV_27 $T=193200 214880 0 0 $X=193010 $Y=214640
X1284 1 2 472 116 ICV_27 $T=212980 182240 0 0 $X=212790 $Y=182000
X1285 1 2 4 476 ICV_27 $T=217580 182240 0 0 $X=217390 $Y=182000
X1286 1 2 183 195 ICV_27 $T=225400 214880 0 0 $X=225210 $Y=214640
X1287 1 2 493 207 ICV_27 $T=253000 204000 0 0 $X=252810 $Y=203760
X1288 1 2 213 214 ICV_27 $T=259440 209440 0 0 $X=259250 $Y=209200
X1289 1 2 505 156 ICV_27 $T=275080 193120 1 0 $X=274890 $Y=190160
X1290 1 2 3 4 ICV_27 $T=337640 193120 0 0 $X=337450 $Y=192880
X1291 1 2 ICV_29 $T=10580 176800 1 0 $X=10390 $Y=173840
X1292 1 2 ICV_29 $T=10580 198560 1 0 $X=10390 $Y=195600
X1293 1 2 ICV_29 $T=10580 209440 1 0 $X=10390 $Y=206480
X1294 1 2 ICV_29 $T=10580 214880 1 0 $X=10390 $Y=211920
X1295 1 2 ICV_29 $T=46000 204000 0 0 $X=45810 $Y=203760
X1296 1 2 ICV_29 $T=65780 187680 1 0 $X=65590 $Y=184720
X1297 1 2 ICV_29 $T=109480 214880 1 0 $X=109290 $Y=211920
X1298 1 2 ICV_29 $T=149500 187680 1 0 $X=149310 $Y=184720
X1299 1 2 ICV_29 $T=164680 209440 0 0 $X=164490 $Y=209200
X1300 1 2 ICV_29 $T=193200 209440 1 0 $X=193010 $Y=206480
X1301 1 2 ICV_29 $T=203780 209440 1 0 $X=203590 $Y=206480
X1302 1 2 ICV_29 $T=213900 193120 0 0 $X=213710 $Y=192880
X1303 1 2 ICV_29 $T=233220 209440 1 0 $X=233030 $Y=206480
X1304 1 2 ICV_29 $T=251160 176800 1 0 $X=250970 $Y=173840
X1305 1 2 ICV_29 $T=261280 193120 1 0 $X=261090 $Y=190160
X1306 1 2 ICV_29 $T=263120 198560 1 0 $X=262930 $Y=195600
X1307 1 2 ICV_29 $T=284280 198560 1 0 $X=284090 $Y=195600
X1308 1 2 ICV_29 $T=290260 176800 1 0 $X=290070 $Y=173840
X1309 1 2 ICV_29 $T=305900 193120 1 0 $X=305710 $Y=190160
X1310 1 2 ICV_29 $T=318780 176800 1 0 $X=318590 $Y=173840
X1311 1 2 ICV_29 $T=318780 182240 1 0 $X=318590 $Y=179280
X1312 1 2 ICV_29 $T=339940 209440 1 0 $X=339750 $Y=206480
X1313 1 2 ICV_32 $T=19780 204000 1 0 $X=19590 $Y=201040
X1314 1 2 ICV_32 $T=47840 182240 1 0 $X=47650 $Y=179280
X1315 1 2 ICV_32 $T=61640 182240 0 0 $X=61450 $Y=182000
X1316 1 2 ICV_32 $T=61640 204000 0 0 $X=61450 $Y=203760
X1317 1 2 ICV_32 $T=103960 187680 1 0 $X=103770 $Y=184720
X1318 1 2 ICV_32 $T=117760 187680 0 0 $X=117570 $Y=187440
X1319 1 2 ICV_32 $T=132020 198560 1 0 $X=131830 $Y=195600
X1320 1 2 ICV_32 $T=160080 209440 1 0 $X=159890 $Y=206480
X1321 1 2 ICV_32 $T=173880 209440 0 0 $X=173690 $Y=209200
X1322 1 2 ICV_32 $T=188140 187680 1 0 $X=187950 $Y=184720
X1323 1 2 ICV_32 $T=188140 204000 1 0 $X=187950 $Y=201040
X1324 1 2 ICV_32 $T=201940 209440 0 0 $X=201750 $Y=209200
X1325 1 2 ICV_32 $T=216200 193120 1 0 $X=216010 $Y=190160
X1326 1 2 ICV_32 $T=244260 193120 1 0 $X=244070 $Y=190160
X1327 1 2 ICV_32 $T=272320 176800 1 0 $X=272130 $Y=173840
X1328 1 2 ICV_32 $T=314180 182240 0 0 $X=313990 $Y=182000
X1329 1 2 ICV_32 $T=328440 209440 1 0 $X=328250 $Y=206480
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186
** N=424 EP=186 IP=3591 FDC=4365
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=150905 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=156345 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=161785 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=167225 $D=191
X4 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 149600 0 0 $X=5330 $Y=149360
X5 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 155040 1 0 $X=5330 $Y=152080
X6 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 155040 0 0 $X=5330 $Y=154800
X7 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 160480 1 0 $X=5330 $Y=157520
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 160480 0 0 $X=5330 $Y=160240
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 165920 1 0 $X=5330 $Y=162960
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 165920 0 0 $X=5330 $Y=165680
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 171360 1 0 $X=5330 $Y=168400
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 171360 0 0 $X=5330 $Y=171120
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 165920 0 0 $X=6710 $Y=165680
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=8740 165920 1 0 $X=8550 $Y=162960
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=34040 160480 0 0 $X=33850 $Y=160240
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=60260 165920 0 0 $X=60070 $Y=165680
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=74520 171360 1 0 $X=74330 $Y=168400
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=78200 171360 1 0 $X=78010 $Y=168400
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=89240 160480 1 0 $X=89050 $Y=157520
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=95220 155040 0 0 $X=95030 $Y=154800
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=106260 160480 1 0 $X=106070 $Y=157520
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=108560 155040 0 0 $X=108370 $Y=154800
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=116380 165920 0 0 $X=116190 $Y=165680
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=129260 160480 0 0 $X=129070 $Y=160240
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=138920 155040 0 0 $X=138730 $Y=154800
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=142600 149600 0 0 $X=142410 $Y=149360
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=142600 171360 0 0 $X=142410 $Y=171120
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 165920 0 0 $X=144250 $Y=165680
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=186760 160480 1 0 $X=186570 $Y=157520
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=207000 165920 1 0 $X=206810 $Y=162960
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228620 171360 0 0 $X=228430 $Y=171120
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 155040 0 0 $X=230270 $Y=154800
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 160480 0 0 $X=230270 $Y=160240
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=232760 165920 1 0 $X=232570 $Y=162960
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=236440 155040 1 0 $X=236250 $Y=152080
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=239200 171360 1 0 $X=239010 $Y=168400
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=251160 149600 0 0 $X=250970 $Y=149360
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=253000 165920 0 0 $X=252810 $Y=165680
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=254840 160480 0 0 $X=254650 $Y=160240
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 165920 1 0 $X=270750 $Y=162960
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=303140 155040 0 0 $X=302950 $Y=154800
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=307280 155040 1 0 $X=307090 $Y=152080
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 155040 0 0 $X=314450 $Y=154800
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 160480 1 0 $X=314450 $Y=157520
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 160480 0 0 $X=314450 $Y=160240
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=316940 155040 1 0 $X=316750 $Y=152080
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=316940 160480 1 0 $X=316750 $Y=157520
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 149600 0 0 $X=340670 $Y=149360
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 149600 1 180 $X=348950 $Y=149360
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 155040 0 180 $X=348950 $Y=152080
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 155040 1 180 $X=348950 $Y=154800
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 160480 0 180 $X=348950 $Y=157520
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 160480 1 180 $X=348950 $Y=160240
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 165920 0 180 $X=348950 $Y=162960
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 165920 1 180 $X=348950 $Y=165680
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 171360 0 180 $X=348950 $Y=168400
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 171360 1 180 $X=348950 $Y=171120
X122 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=12420 171360 0 0 $X=12230 $Y=171120
X123 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 155040 1 0 $X=15910 $Y=152080
X124 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=28980 149600 0 0 $X=28790 $Y=149360
X125 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39560 149600 0 0 $X=39370 $Y=149360
X126 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 171360 1 0 $X=43970 $Y=168400
X127 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44620 155040 0 0 $X=44430 $Y=154800
X128 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=46460 171360 0 0 $X=46270 $Y=171120
X129 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=49220 155040 0 0 $X=49030 $Y=154800
X130 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=56580 165920 0 0 $X=56390 $Y=165680
X131 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57500 149600 0 0 $X=57310 $Y=149360
X132 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57500 160480 1 0 $X=57310 $Y=157520
X133 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 171360 0 0 $X=57770 $Y=171120
X134 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=65780 155040 0 0 $X=65590 $Y=154800
X135 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=70840 149600 0 0 $X=70650 $Y=149360
X136 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 155040 1 0 $X=72030 $Y=152080
X137 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 160480 1 0 $X=72030 $Y=157520
X138 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 165920 1 0 $X=72030 $Y=162960
X139 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 165920 1 0 $X=76170 $Y=162960
X140 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 171360 1 0 $X=89970 $Y=168400
X141 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 160480 1 0 $X=100090 $Y=157520
X142 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=107640 149600 0 0 $X=107450 $Y=149360
X143 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=108560 171360 0 0 $X=108370 $Y=171120
X144 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=113160 171360 0 0 $X=112970 $Y=171120
X145 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=125580 165920 1 0 $X=125390 $Y=162960
X146 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=127420 160480 1 0 $X=127230 $Y=157520
X147 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=127880 155040 1 0 $X=127690 $Y=152080
X148 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 155040 1 0 $X=132290 $Y=152080
X149 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=154560 171360 1 0 $X=154370 $Y=168400
X150 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=162840 171360 1 0 $X=162650 $Y=168400
X151 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=171120 165920 1 0 $X=170930 $Y=162960
X152 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178020 160480 1 0 $X=177830 $Y=157520
X153 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178020 171360 1 0 $X=177830 $Y=168400
X154 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183080 160480 1 0 $X=182890 $Y=157520
X155 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194120 165920 1 0 $X=193930 $Y=162960
X156 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=197340 165920 0 0 $X=197150 $Y=165680
X157 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=202400 160480 0 0 $X=202210 $Y=160240
X158 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=203780 171360 1 0 $X=203590 $Y=168400
X159 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=207000 160480 1 0 $X=206810 $Y=157520
X160 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=210680 171360 1 0 $X=210490 $Y=168400
X161 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212060 155040 0 0 $X=211870 $Y=154800
X162 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 165920 1 0 $X=212330 $Y=162960
X163 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=213440 149600 0 0 $X=213250 $Y=149360
X164 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=222180 155040 1 0 $X=221990 $Y=152080
X165 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=228620 171360 1 0 $X=228430 $Y=168400
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=232300 171360 0 0 $X=232110 $Y=171120
X167 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239660 160480 1 0 $X=239470 $Y=157520
X168 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 165920 1 0 $X=240390 $Y=162960
X169 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=242880 160480 0 0 $X=242690 $Y=160240
X170 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249320 165920 0 0 $X=249130 $Y=165680
X171 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=261740 155040 1 0 $X=261550 $Y=152080
X172 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=262200 165920 1 0 $X=262010 $Y=162960
X173 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267260 165920 1 0 $X=267070 $Y=162960
X174 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 155040 1 0 $X=268450 $Y=152080
X175 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 160480 1 0 $X=268450 $Y=157520
X176 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 171360 1 0 $X=268450 $Y=168400
X177 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=270940 149600 0 0 $X=270750 $Y=149360
X178 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=270940 165920 0 0 $X=270750 $Y=165680
X179 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 171360 1 0 $X=272590 $Y=168400
X180 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=277840 149600 0 0 $X=277650 $Y=149360
X181 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=294860 155040 1 0 $X=294670 $Y=152080
X182 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 171360 1 0 $X=296510 $Y=168400
X183 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 171360 1 0 $X=300650 $Y=168400
X184 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 171360 0 0 $X=300650 $Y=171120
X185 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=321540 165920 0 0 $X=321350 $Y=165680
X186 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 155040 1 0 $X=324570 $Y=152080
X187 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 160480 1 0 $X=324570 $Y=157520
X188 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=338560 171360 0 0 $X=338370 $Y=171120
X189 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 155040 1 0 $X=345270 $Y=152080
X190 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 160480 1 0 $X=345270 $Y=157520
X191 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 165920 1 0 $X=345270 $Y=162960
X192 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 171360 1 0 $X=345270 $Y=168400
X193 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 171360 0 0 $X=6710 $Y=171120
X194 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=10580 155040 1 0 $X=10390 $Y=152080
X195 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=29440 171360 1 0 $X=29250 $Y=168400
X196 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=31740 160480 1 0 $X=31550 $Y=157520
X197 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=33580 165920 1 0 $X=33390 $Y=162960
X198 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=39100 155040 0 0 $X=38910 $Y=154800
X199 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40020 160480 1 0 $X=39830 $Y=157520
X200 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55660 165920 1 0 $X=55470 $Y=162960
X201 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=59340 155040 1 0 $X=59150 $Y=152080
X202 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=59800 171360 1 0 $X=59610 $Y=168400
X203 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=70380 165920 0 0 $X=70190 $Y=165680
X204 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81420 155040 0 0 $X=81230 $Y=154800
X205 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=89700 155040 1 0 $X=89510 $Y=152080
X206 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=118680 171360 1 0 $X=118490 $Y=168400
X207 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=120060 165920 1 0 $X=119870 $Y=162960
X208 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=121900 160480 1 0 $X=121710 $Y=157520
X209 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 155040 0 0 $X=125390 $Y=154800
X210 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=129720 149600 0 0 $X=129530 $Y=149360
X211 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=162380 149600 0 0 $X=162190 $Y=149360
X212 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=169280 160480 1 0 $X=169090 $Y=157520
X213 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=180780 149600 0 0 $X=180590 $Y=149360
X214 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=195500 149600 0 0 $X=195310 $Y=149360
X215 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=200100 165920 1 0 $X=199910 $Y=162960
X216 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210680 155040 1 0 $X=210490 $Y=152080
X217 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=223100 160480 1 0 $X=222910 $Y=157520
X218 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=225860 165920 1 0 $X=225670 $Y=162960
X219 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=230000 155040 1 0 $X=229810 $Y=152080
X220 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=233680 171360 1 0 $X=233490 $Y=168400
X221 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=238740 149600 0 0 $X=238550 $Y=149360
X222 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=263120 160480 1 0 $X=262930 $Y=157520
X223 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=275540 155040 0 0 $X=275350 $Y=154800
X224 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=295320 171360 0 0 $X=295130 $Y=171120
X225 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=297620 155040 0 0 $X=297430 $Y=154800
X226 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322460 171360 1 0 $X=322270 $Y=168400
X227 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=325680 171360 0 0 $X=325490 $Y=171120
X228 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=335340 149600 0 0 $X=335150 $Y=149360
X229 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=339940 155040 1 0 $X=339750 $Y=152080
X230 1 2 ICV_2 $T=33580 149600 0 0 $X=33390 $Y=149360
X231 1 2 ICV_2 $T=33580 165920 0 0 $X=33390 $Y=165680
X232 1 2 ICV_2 $T=61640 149600 0 0 $X=61450 $Y=149360
X233 1 2 ICV_2 $T=89700 171360 0 0 $X=89510 $Y=171120
X234 1 2 ICV_2 $T=103960 155040 1 0 $X=103770 $Y=152080
X235 1 2 ICV_2 $T=117760 171360 0 0 $X=117570 $Y=171120
X236 1 2 ICV_2 $T=188140 165920 1 0 $X=187950 $Y=162960
X237 1 2 ICV_2 $T=216200 155040 1 0 $X=216010 $Y=152080
X238 1 2 ICV_2 $T=230000 149600 0 0 $X=229810 $Y=149360
X239 1 2 ICV_2 $T=244260 160480 1 0 $X=244070 $Y=157520
X240 1 2 ICV_2 $T=244260 165920 1 0 $X=244070 $Y=162960
X241 1 2 ICV_2 $T=272320 165920 1 0 $X=272130 $Y=162960
X242 1 2 ICV_2 $T=300380 160480 1 0 $X=300190 $Y=157520
X243 1 2 ICV_2 $T=328440 160480 1 0 $X=328250 $Y=157520
X244 1 2 ICV_2 $T=328440 165920 1 0 $X=328250 $Y=162960
X245 1 2 ICV_2 $T=328440 171360 1 0 $X=328250 $Y=168400
X246 1 2 ICV_2 $T=342240 149600 0 0 $X=342050 $Y=149360
X247 1 2 ICV_2 $T=342240 155040 0 0 $X=342050 $Y=154800
X248 1 2 ICV_2 $T=342240 160480 0 0 $X=342050 $Y=160240
X249 1 2 ICV_2 $T=342240 165920 0 0 $X=342050 $Y=165680
X250 1 2 ICV_2 $T=342240 171360 0 0 $X=342050 $Y=171120
X251 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 171360 1 0 $X=17750 $Y=168400
X252 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 160480 0 0 $X=18210 $Y=160240
X253 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=20700 165920 0 0 $X=20510 $Y=165680
X254 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 171360 0 0 $X=33850 $Y=171120
X255 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 155040 1 0 $X=45810 $Y=152080
X256 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 165920 0 0 $X=61910 $Y=165680
X257 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 160480 1 0 $X=76170 $Y=157520
X258 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=81880 155040 1 0 $X=81690 $Y=152080
X259 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=82800 165920 1 0 $X=82610 $Y=162960
X260 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=93380 160480 1 0 $X=93190 $Y=157520
X261 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=93840 149600 0 0 $X=93650 $Y=149360
X262 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 160480 0 0 $X=101930 $Y=160240
X263 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=103960 155040 0 0 $X=103770 $Y=154800
X264 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=112700 155040 1 0 $X=112510 $Y=152080
X265 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=124200 171360 1 0 $X=124010 $Y=168400
X266 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=127880 171360 0 0 $X=127690 $Y=171120
X267 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=141680 155040 0 0 $X=141490 $Y=154800
X268 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143060 171360 1 0 $X=142870 $Y=168400
X269 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=146280 160480 0 0 $X=146090 $Y=160240
X270 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 160480 1 0 $X=160350 $Y=157520
X271 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=165600 165920 0 0 $X=165410 $Y=165680
X272 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=167900 149600 0 0 $X=167710 $Y=149360
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174340 155040 0 0 $X=174150 $Y=154800
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174340 171360 0 0 $X=174150 $Y=171120
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174800 160480 1 0 $X=174610 $Y=157520
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=179400 165920 0 0 $X=179210 $Y=165680
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188140 165920 0 0 $X=187950 $Y=165680
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188600 160480 1 0 $X=188410 $Y=157520
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 160480 1 0 $X=214170 $Y=157520
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 171360 1 0 $X=216470 $Y=168400
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=220340 171360 0 0 $X=220150 $Y=171120
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 165920 0 0 $X=242230 $Y=165680
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=250240 160480 0 0 $X=250050 $Y=160240
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 149600 0 0 $X=258330 $Y=149360
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 171360 1 0 $X=258330 $Y=168400
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 171360 0 0 $X=258330 $Y=171120
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=272320 160480 0 0 $X=272130 $Y=160240
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=281060 165920 1 0 $X=280870 $Y=162960
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=283820 155040 1 0 $X=283630 $Y=152080
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286580 165920 0 0 $X=286390 $Y=165680
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 160480 1 0 $X=298350 $Y=157520
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=301300 160480 0 0 $X=301110 $Y=160240
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=332580 155040 0 0 $X=332390 $Y=154800
X294 1 4 sky130_fd_sc_hd__diode_2 $T=7820 165920 1 0 $X=7630 $Y=162960
X295 1 4 sky130_fd_sc_hd__diode_2 $T=8280 165920 0 0 $X=8090 $Y=165680
X296 1 4 sky130_fd_sc_hd__diode_2 $T=19320 155040 0 0 $X=19130 $Y=154800
X297 1 14 sky130_fd_sc_hd__diode_2 $T=21160 171360 1 0 $X=20970 $Y=168400
X298 1 16 sky130_fd_sc_hd__diode_2 $T=23920 160480 0 0 $X=23730 $Y=160240
X299 1 322 sky130_fd_sc_hd__diode_2 $T=26220 165920 1 0 $X=26030 $Y=162960
X300 1 329 sky130_fd_sc_hd__diode_2 $T=48300 155040 0 0 $X=48110 $Y=154800
X301 1 33 sky130_fd_sc_hd__diode_2 $T=64400 165920 0 0 $X=64210 $Y=165680
X302 1 34 sky130_fd_sc_hd__diode_2 $T=64860 171360 0 0 $X=64670 $Y=171120
X303 1 332 sky130_fd_sc_hd__diode_2 $T=66240 165920 1 0 $X=66050 $Y=162960
X304 1 37 sky130_fd_sc_hd__diode_2 $T=69920 155040 0 0 $X=69730 $Y=154800
X305 1 39 sky130_fd_sc_hd__diode_2 $T=72680 171360 0 0 $X=72490 $Y=171120
X306 1 334 sky130_fd_sc_hd__diode_2 $T=77280 171360 1 0 $X=77090 $Y=168400
X307 1 52 sky130_fd_sc_hd__diode_2 $T=93840 160480 0 0 $X=93650 $Y=160240
X308 1 54 sky130_fd_sc_hd__diode_2 $T=96600 155040 0 0 $X=96410 $Y=154800
X309 1 343 sky130_fd_sc_hd__diode_2 $T=99360 160480 1 0 $X=99170 $Y=157520
X310 1 57 sky130_fd_sc_hd__diode_2 $T=101660 149600 0 0 $X=101470 $Y=149360
X311 1 338 sky130_fd_sc_hd__diode_2 $T=102580 171360 0 0 $X=102390 $Y=171120
X312 1 49 sky130_fd_sc_hd__diode_2 $T=103500 165920 0 0 $X=103310 $Y=165680
X313 1 347 sky130_fd_sc_hd__diode_2 $T=105340 160480 1 0 $X=105150 $Y=157520
X314 1 345 sky130_fd_sc_hd__diode_2 $T=108100 160480 0 0 $X=107910 $Y=160240
X315 1 349 sky130_fd_sc_hd__diode_2 $T=110400 171360 1 0 $X=110210 $Y=168400
X316 1 351 sky130_fd_sc_hd__diode_2 $T=112240 171360 0 0 $X=112050 $Y=171120
X317 1 62 sky130_fd_sc_hd__diode_2 $T=112700 165920 1 0 $X=112510 $Y=162960
X318 1 353 sky130_fd_sc_hd__diode_2 $T=115460 165920 0 0 $X=115270 $Y=165680
X319 1 44 sky130_fd_sc_hd__diode_2 $T=124660 171360 0 0 $X=124470 $Y=171120
X320 1 357 sky130_fd_sc_hd__diode_2 $T=135700 149600 0 0 $X=135510 $Y=149360
X321 1 75 sky130_fd_sc_hd__diode_2 $T=135700 171360 1 0 $X=135510 $Y=168400
X322 1 358 sky130_fd_sc_hd__diode_2 $T=138000 155040 0 0 $X=137810 $Y=154800
X323 1 70 sky130_fd_sc_hd__diode_2 $T=149500 165920 0 0 $X=149310 $Y=165680
X324 1 87 sky130_fd_sc_hd__diode_2 $T=149960 171360 0 0 $X=149770 $Y=171120
X325 1 89 sky130_fd_sc_hd__diode_2 $T=154560 155040 0 0 $X=154370 $Y=154800
X326 1 88 sky130_fd_sc_hd__diode_2 $T=162840 160480 0 0 $X=162650 $Y=160240
X327 1 106 sky130_fd_sc_hd__diode_2 $T=189520 149600 0 0 $X=189330 $Y=149360
X328 1 79 sky130_fd_sc_hd__diode_2 $T=190440 165920 0 0 $X=190250 $Y=165680
X329 1 368 sky130_fd_sc_hd__diode_2 $T=206080 165920 1 0 $X=205890 $Y=162960
X330 1 353 sky130_fd_sc_hd__diode_2 $T=209760 160480 0 0 $X=209570 $Y=160240
X331 1 66 sky130_fd_sc_hd__diode_2 $T=209760 171360 1 0 $X=209570 $Y=168400
X332 1 131 sky130_fd_sc_hd__diode_2 $T=222640 165920 1 0 $X=222450 $Y=162960
X333 1 138 sky130_fd_sc_hd__diode_2 $T=231380 165920 0 0 $X=231190 $Y=165680
X334 1 137 sky130_fd_sc_hd__diode_2 $T=231380 171360 0 0 $X=231190 $Y=171120
X335 1 139 sky130_fd_sc_hd__diode_2 $T=231840 155040 0 0 $X=231650 $Y=154800
X336 1 375 sky130_fd_sc_hd__diode_2 $T=231840 165920 1 0 $X=231650 $Y=162960
X337 1 376 sky130_fd_sc_hd__diode_2 $T=235520 155040 1 0 $X=235330 $Y=152080
X338 1 138 sky130_fd_sc_hd__diode_2 $T=239200 165920 0 0 $X=239010 $Y=165680
X339 1 375 sky130_fd_sc_hd__diode_2 $T=241960 160480 0 0 $X=241770 $Y=160240
X340 1 138 sky130_fd_sc_hd__diode_2 $T=247020 160480 0 0 $X=246830 $Y=160240
X341 1 141 sky130_fd_sc_hd__diode_2 $T=248400 165920 0 0 $X=248210 $Y=165680
X342 1 379 sky130_fd_sc_hd__diode_2 $T=251160 160480 1 0 $X=250970 $Y=157520
X343 1 380 sky130_fd_sc_hd__diode_2 $T=261280 165920 1 0 $X=261090 $Y=162960
X344 1 382 sky130_fd_sc_hd__diode_2 $T=264500 155040 0 0 $X=264310 $Y=154800
X345 1 64 sky130_fd_sc_hd__diode_2 $T=267720 155040 1 0 $X=267530 $Y=152080
X346 1 145 sky130_fd_sc_hd__diode_2 $T=276920 149600 0 0 $X=276730 $Y=149360
X347 1 389 sky130_fd_sc_hd__diode_2 $T=285200 160480 1 0 $X=285010 $Y=157520
X348 1 149 sky130_fd_sc_hd__diode_2 $T=287500 149600 0 0 $X=287310 $Y=149360
X349 1 147 sky130_fd_sc_hd__diode_2 $T=288880 165920 0 0 $X=288690 $Y=165680
X350 1 170 sky130_fd_sc_hd__diode_2 $T=304520 155040 0 0 $X=304330 $Y=154800
X351 1 172 sky130_fd_sc_hd__diode_2 $T=304520 171360 0 0 $X=304330 $Y=171120
X352 1 395 sky130_fd_sc_hd__diode_2 $T=306360 155040 1 0 $X=306170 $Y=152080
X353 1 175 sky130_fd_sc_hd__diode_2 $T=307280 160480 1 0 $X=307090 $Y=157520
X354 1 171 sky130_fd_sc_hd__diode_2 $T=308660 155040 1 0 $X=308470 $Y=152080
X355 1 170 sky130_fd_sc_hd__diode_2 $T=316020 160480 1 0 $X=315830 $Y=157520
X356 1 402 sky130_fd_sc_hd__diode_2 $T=326140 165920 0 0 $X=325950 $Y=165680
X357 1 183 sky130_fd_sc_hd__diode_2 $T=337640 171360 0 0 $X=337450 $Y=171120
X358 1 2 323 ICV_4 $T=30360 165920 0 0 $X=30170 $Y=165680
X359 1 2 18 ICV_4 $T=30820 160480 0 0 $X=30630 $Y=160240
X360 1 2 17 ICV_4 $T=30820 171360 0 0 $X=30630 $Y=171120
X361 1 2 28 ICV_4 $T=51060 171360 0 0 $X=50870 $Y=171120
X362 1 2 325 ICV_4 $T=52900 160480 1 0 $X=52710 $Y=157520
X363 1 2 46 ICV_4 $T=81880 171360 1 0 $X=81690 $Y=168400
X364 1 2 48 ICV_4 $T=86480 149600 0 0 $X=86290 $Y=149360
X365 1 2 49 ICV_4 $T=86480 165920 0 0 $X=86290 $Y=165680
X366 1 2 52 ICV_4 $T=91080 160480 0 0 $X=90890 $Y=160240
X367 1 2 55 ICV_4 $T=100280 165920 0 0 $X=100090 $Y=165680
X368 1 2 53 ICV_4 $T=100740 155040 1 0 $X=100550 $Y=152080
X369 1 2 65 ICV_4 $T=115000 160480 0 0 $X=114810 $Y=160240
X370 1 2 55 ICV_4 $T=133860 165920 0 0 $X=133670 $Y=165680
X371 1 2 70 ICV_4 $T=143060 160480 0 0 $X=142870 $Y=160240
X372 1 2 359 ICV_4 $T=145820 165920 1 0 $X=145630 $Y=162960
X373 1 2 75 ICV_4 $T=147200 171360 0 0 $X=147010 $Y=171120
X374 1 2 80 ICV_4 $T=147660 160480 1 0 $X=147470 $Y=157520
X375 1 2 86 ICV_4 $T=148580 171360 1 0 $X=148390 $Y=168400
X376 1 2 362 ICV_4 $T=155020 165920 1 0 $X=154830 $Y=162960
X377 1 2 55 ICV_4 $T=161460 165920 1 0 $X=161270 $Y=162960
X378 1 2 92 ICV_4 $T=171120 160480 0 0 $X=170930 $Y=160240
X379 1 2 89 ICV_4 $T=182620 155040 0 0 $X=182430 $Y=154800
X380 1 2 111 ICV_4 $T=193660 155040 0 0 $X=193470 $Y=154800
X381 1 2 118 ICV_4 $T=198720 160480 0 0 $X=198530 $Y=160240
X382 1 2 85 ICV_4 $T=199180 155040 0 0 $X=198990 $Y=154800
X383 1 2 120 ICV_4 $T=199180 171360 0 0 $X=198990 $Y=171120
X384 1 2 129 ICV_4 $T=226780 165920 0 0 $X=226590 $Y=165680
X385 1 2 381 ICV_4 $T=253000 155040 1 0 $X=252810 $Y=152080
X386 1 2 351 ICV_4 $T=254840 155040 0 0 $X=254650 $Y=154800
X387 1 2 65 ICV_4 $T=261740 165920 0 0 $X=261550 $Y=165680
X388 1 2 166 ICV_4 $T=303600 160480 0 0 $X=303410 $Y=160240
X389 1 2 394 ICV_4 $T=305900 165920 1 0 $X=305710 $Y=162960
X390 1 2 101 ICV_4 $T=311420 155040 0 0 $X=311230 $Y=154800
X391 1 2 170 ICV_4 $T=311420 165920 0 0 $X=311230 $Y=165680
X392 1 2 4 ICV_4 $T=311420 171360 0 0 $X=311230 $Y=171120
X393 1 2 397 ICV_4 $T=315560 165920 0 0 $X=315370 $Y=165680
X394 1 2 401 ICV_4 $T=325220 165920 1 0 $X=325030 $Y=162960
X395 1 2 402 ICV_4 $T=339020 160480 0 0 $X=338830 $Y=160240
X396 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 165920 1 0 $X=16370 $Y=162960
X397 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=25300 155040 0 0 $X=25110 $Y=154800
X398 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58880 155040 0 0 $X=58690 $Y=154800
X399 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=62100 171360 0 0 $X=61910 $Y=171120
X400 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=64860 155040 1 0 $X=64670 $Y=152080
X401 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=65320 171360 1 0 $X=65130 $Y=168400
X402 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=75900 155040 0 0 $X=75710 $Y=154800
X403 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=76360 155040 1 0 $X=76170 $Y=152080
X404 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=87400 165920 1 0 $X=87210 $Y=162960
X405 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=98440 149600 0 0 $X=98250 $Y=149360
X406 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=98900 171360 1 0 $X=98710 $Y=168400
X407 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=131100 155040 0 0 $X=130910 $Y=154800
X408 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157320 160480 1 0 $X=157130 $Y=157520
X409 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=167440 171360 0 0 $X=167250 $Y=171120
X410 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=171580 155040 1 0 $X=171390 $Y=152080
X411 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=186300 149600 0 0 $X=186110 $Y=149360
X412 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 155040 0 0 $X=202210 $Y=154800
X413 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 171360 0 0 $X=202210 $Y=171120
X414 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202860 160480 1 0 $X=202670 $Y=157520
X415 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=225400 160480 0 0 $X=225210 $Y=160240
X416 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 155040 0 0 $X=226590 $Y=154800
X417 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=228620 160480 1 0 $X=228430 $Y=157520
X418 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=249780 155040 1 0 $X=249590 $Y=152080
X419 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=251160 171360 1 0 $X=250970 $Y=168400
X420 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=281060 155040 0 0 $X=280870 $Y=154800
X421 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297160 165920 1 0 $X=296970 $Y=162960
X422 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 165920 1 0 $X=300650 $Y=162960
X423 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=303140 155040 1 0 $X=302950 $Y=152080
X424 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=312800 171360 1 0 $X=312610 $Y=168400
X425 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 149600 0 0 $X=314450 $Y=149360
X426 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331200 171360 0 0 $X=331010 $Y=171120
X427 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=332120 165920 0 0 $X=331930 $Y=165680
X428 1 2 13 ICV_5 $T=28060 155040 0 0 $X=27870 $Y=154800
X429 1 2 4 ICV_5 $T=35880 171360 1 0 $X=35690 $Y=168400
X430 1 2 27 ICV_5 $T=55660 160480 0 0 $X=55470 $Y=160240
X431 1 2 330 ICV_5 $T=62100 165920 1 0 $X=61910 $Y=162960
X432 1 2 36 ICV_5 $T=74520 160480 0 0 $X=74330 $Y=160240
X433 1 2 47 ICV_5 $T=85560 171360 0 0 $X=85370 $Y=171120
X434 1 2 344 ICV_5 $T=97980 165920 1 0 $X=97790 $Y=162960
X435 1 2 44 ICV_5 $T=98900 171360 0 0 $X=98710 $Y=171120
X436 1 2 83 ICV_5 $T=152260 155040 1 0 $X=152070 $Y=152080
X437 1 2 88 ICV_5 $T=156400 155040 1 0 $X=156210 $Y=152080
X438 1 2 87 ICV_5 $T=175260 160480 0 0 $X=175070 $Y=160240
X439 1 2 102 ICV_5 $T=176640 155040 0 0 $X=176450 $Y=154800
X440 1 2 107 ICV_5 $T=184000 171360 1 0 $X=183810 $Y=168400
X441 1 2 134 ICV_5 $T=225860 149600 0 0 $X=225670 $Y=149360
X442 1 2 132 ICV_5 $T=235520 165920 0 0 $X=235330 $Y=165680
X443 1 2 378 ICV_5 $T=240120 155040 1 0 $X=239930 $Y=152080
X444 1 2 130 ICV_5 $T=240580 171360 1 0 $X=240390 $Y=168400
X445 1 2 4 ICV_5 $T=260820 171360 1 0 $X=260630 $Y=168400
X446 1 2 127 ICV_5 $T=268640 155040 0 0 $X=268450 $Y=154800
X447 1 2 159 ICV_5 $T=304980 171360 1 0 $X=304790 $Y=168400
X448 1 2 120 ICV_5 $T=338560 155040 0 0 $X=338370 $Y=154800
X449 1 2 182 ICV_5 $T=338560 165920 0 0 $X=338370 $Y=165680
X450 1 3 4 ICV_7 $T=7820 155040 1 0 $X=7630 $Y=152080
X451 1 3 5 ICV_7 $T=7820 160480 1 0 $X=7630 $Y=157520
X452 1 7 10 ICV_7 $T=17020 171360 0 0 $X=16830 $Y=171120
X453 1 11 321 ICV_7 $T=20240 160480 0 0 $X=20050 $Y=160240
X454 1 13 15 ICV_7 $T=20700 171360 0 0 $X=20510 $Y=171120
X455 1 320 12 ICV_7 $T=21160 155040 1 0 $X=20970 $Y=152080
X456 1 10 17 ICV_7 $T=23000 165920 0 0 $X=22810 $Y=165680
X457 1 7 321 ICV_7 $T=26680 165920 0 0 $X=26490 $Y=165680
X458 1 324 21 ICV_7 $T=35420 160480 0 0 $X=35230 $Y=160240
X459 1 16 326 ICV_7 $T=40020 165920 0 0 $X=39830 $Y=165680
X460 1 23 4 ICV_7 $T=43240 149600 0 0 $X=43050 $Y=149360
X461 1 327 4 ICV_7 $T=43700 165920 0 0 $X=43510 $Y=165680
X462 1 21 22 ICV_7 $T=49220 160480 1 0 $X=49030 $Y=157520
X463 1 26 27 ICV_7 $T=53820 165920 0 0 $X=53630 $Y=165680
X464 1 31 29 ICV_7 $T=56120 155040 0 0 $X=55930 $Y=154800
X465 1 4 331 ICV_7 $T=63020 155040 0 0 $X=62830 $Y=154800
X466 1 33 333 ICV_7 $T=68080 149600 0 0 $X=67890 $Y=149360
X467 1 35 38 ICV_7 $T=69000 171360 0 0 $X=68810 $Y=171120
X468 1 335 41 ICV_7 $T=75440 149600 0 0 $X=75250 $Y=149360
X469 1 40 42 ICV_7 $T=76360 165920 0 0 $X=76170 $Y=165680
X470 1 336 338 ICV_7 $T=78200 160480 0 0 $X=78010 $Y=160240
X471 1 4 337 ICV_7 $T=78660 155040 0 0 $X=78470 $Y=154800
X472 1 43 339 ICV_7 $T=79120 155040 1 0 $X=78930 $Y=152080
X473 1 334 44 ICV_7 $T=80040 165920 1 0 $X=79850 $Y=162960
X474 1 39 38 ICV_7 $T=81880 171360 0 0 $X=81690 $Y=171120
X475 1 40 46 ICV_7 $T=84640 165920 1 0 $X=84450 $Y=162960
X476 1 51 341 ICV_7 $T=90620 160480 1 0 $X=90430 $Y=157520
X477 1 40 335 ICV_7 $T=91080 149600 0 0 $X=90890 $Y=149360
X478 1 53 340 ICV_7 $T=93840 171360 1 0 $X=93650 $Y=168400
X479 1 338 342 ICV_7 $T=95680 149600 0 0 $X=95490 $Y=149360
X480 1 51 343 ICV_7 $T=95680 160480 1 0 $X=95490 $Y=157520
X481 1 52 51 ICV_7 $T=104420 160480 0 0 $X=104230 $Y=160240
X482 1 348 4 ICV_7 $T=105800 155040 0 0 $X=105610 $Y=154800
X483 1 338 350 ICV_7 $T=109940 155040 1 0 $X=109750 $Y=152080
X484 1 338 53 ICV_7 $T=111780 165920 0 0 $X=111590 $Y=165680
X485 1 60 64 ICV_7 $T=112240 149600 0 0 $X=112050 $Y=149360
X486 1 351 60 ICV_7 $T=119140 160480 1 0 $X=118950 $Y=157520
X487 1 53 62 ICV_7 $T=119140 160480 0 0 $X=118950 $Y=160240
X488 1 67 68 ICV_7 $T=126500 171360 1 0 $X=126310 $Y=168400
X489 1 354 70 ICV_7 $T=127880 165920 0 0 $X=127690 $Y=165680
X490 1 71 73 ICV_7 $T=129720 171360 0 0 $X=129530 $Y=171120
X491 1 355 55 ICV_7 $T=130640 160480 0 0 $X=130450 $Y=160240
X492 1 74 4 ICV_7 $T=134320 155040 0 0 $X=134130 $Y=154800
X493 1 29 31 ICV_7 $T=134320 160480 0 0 $X=134130 $Y=160240
X494 1 4 77 ICV_7 $T=139840 149600 0 0 $X=139650 $Y=149360
X495 1 80 72 ICV_7 $T=139840 171360 0 0 $X=139650 $Y=171120
X496 1 79 71 ICV_7 $T=141680 165920 0 0 $X=141490 $Y=165680
X497 1 67 80 ICV_7 $T=144900 171360 1 0 $X=144710 $Y=168400
X498 1 360 361 ICV_7 $T=148580 155040 1 0 $X=148390 $Y=152080
X499 1 85 88 ICV_7 $T=148580 160480 0 0 $X=148390 $Y=160240
X500 1 82 88 ICV_7 $T=151800 171360 1 0 $X=151610 $Y=168400
X501 1 91 94 ICV_7 $T=158240 171360 0 0 $X=158050 $Y=171120
X502 1 364 365 ICV_7 $T=159160 160480 0 0 $X=158970 $Y=160240
X503 1 95 90 ICV_7 $T=162840 160480 1 0 $X=162650 $Y=157520
X504 1 365 366 ICV_7 $T=166520 160480 1 0 $X=166330 $Y=157520
X505 1 4 363 ICV_7 $T=167440 165920 0 0 $X=167250 $Y=165680
X506 1 96 25 ICV_7 $T=170200 149600 0 0 $X=170010 $Y=149360
X507 1 97 99 ICV_7 $T=170200 171360 0 0 $X=170010 $Y=171120
X508 1 108 102 ICV_7 $T=187680 155040 0 0 $X=187490 $Y=154800
X509 1 109 106 ICV_7 $T=189520 171360 1 0 $X=189330 $Y=168400
X510 1 4 367 ICV_7 $T=194580 165920 0 0 $X=194390 $Y=165680
X511 1 116 113 ICV_7 $T=195500 171360 0 0 $X=195310 $Y=171120
X512 1 122 369 ICV_7 $T=206080 160480 0 0 $X=205890 $Y=160240
X513 1 351 372 ICV_7 $T=211600 160480 1 0 $X=211410 $Y=157520
X514 1 371 125 ICV_7 $T=212520 171360 0 0 $X=212330 $Y=171120
X515 1 127 123 ICV_7 $T=216660 155040 0 0 $X=216470 $Y=154800
X516 1 129 123 ICV_7 $T=218500 171360 1 0 $X=218310 $Y=168400
X517 1 125 370 ICV_7 $T=218960 160480 0 0 $X=218770 $Y=160240
X518 1 373 133 ICV_7 $T=222180 171360 0 0 $X=221990 $Y=171120
X519 1 130 132 ICV_7 $T=222640 160480 0 0 $X=222450 $Y=160240
X520 1 131 130 ICV_7 $T=225860 171360 0 0 $X=225670 $Y=171120
X521 1 89 374 ICV_7 $T=231840 160480 1 0 $X=231650 $Y=157520
X522 1 132 4 ICV_7 $T=235980 155040 0 0 $X=235790 $Y=154800
X523 1 377 131 ICV_7 $T=236900 171360 0 0 $X=236710 $Y=171120
X524 1 131 130 ICV_7 $T=238280 160480 0 0 $X=238090 $Y=160240
X525 1 79 123 ICV_7 $T=244720 165920 0 0 $X=244530 $Y=165680
X526 1 73 143 ICV_7 $T=247940 171360 0 0 $X=247750 $Y=171120
X527 1 144 353 ICV_7 $T=251160 155040 0 0 $X=250970 $Y=154800
X528 1 351 353 ICV_7 $T=252080 160480 0 0 $X=251890 $Y=160240
X529 1 144 145 ICV_7 $T=252540 149600 0 0 $X=252350 $Y=149360
X530 1 125 383 ICV_7 $T=254380 165920 0 0 $X=254190 $Y=165680
X531 1 125 123 ICV_7 $T=260360 160480 1 0 $X=260170 $Y=157520
X532 1 4 385 ICV_7 $T=272780 155040 0 0 $X=272590 $Y=154800
X533 1 386 154 ICV_7 $T=274620 160480 0 0 $X=274430 $Y=160240
X534 1 387 4 ICV_7 $T=274620 165920 0 0 $X=274430 $Y=165680
X535 1 154 388 ICV_7 $T=278300 165920 1 0 $X=278110 $Y=162960
X536 1 155 159 ICV_7 $T=282440 149600 0 0 $X=282250 $Y=149360
X537 1 157 390 ICV_7 $T=283360 165920 1 0 $X=283170 $Y=162960
X538 1 161 162 ICV_7 $T=285660 155040 1 0 $X=285470 $Y=152080
X539 1 157 159 ICV_7 $T=287500 155040 0 0 $X=287310 $Y=154800
X540 1 165 391 ICV_7 $T=292560 171360 0 0 $X=292370 $Y=171120
X541 1 150 159 ICV_7 $T=294400 165920 1 0 $X=294210 $Y=162960
X542 1 169 396 ICV_7 $T=304980 149600 0 0 $X=304790 $Y=149360
X543 1 174 176 ICV_7 $T=306820 160480 0 0 $X=306630 $Y=160240
X544 1 175 176 ICV_7 $T=308660 149600 0 0 $X=308470 $Y=149360
X545 1 394 393 ICV_7 $T=310500 160480 0 0 $X=310310 $Y=160240
X546 1 176 103 ICV_7 $T=316020 155040 0 0 $X=315830 $Y=154800
X547 1 178 176 ICV_7 $T=317400 149600 0 0 $X=317210 $Y=149360
X548 1 174 400 ICV_7 $T=318320 155040 1 0 $X=318130 $Y=152080
X549 1 400 171 ICV_7 $T=318780 165920 0 0 $X=318590 $Y=165680
X550 1 171 178 ICV_7 $T=322000 155040 1 0 $X=321810 $Y=152080
X551 1 3 4 ICV_7 $T=333960 171360 0 0 $X=333770 $Y=171120
X552 1 3 4 ICV_7 $T=334880 155040 0 0 $X=334690 $Y=154800
X553 1 3 4 ICV_7 $T=334880 165920 0 0 $X=334690 $Y=165680
X554 1 3 4 ICV_7 $T=335340 160480 0 0 $X=335150 $Y=160240
X555 1 2 3 5 4 2 8 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 155040 0 0 $X=7630 $Y=154800
X556 1 2 3 6 4 2 9 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 160480 0 0 $X=7630 $Y=160240
X557 1 2 403 318 4 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=10120 165920 0 0 $X=9930 $Y=165680
X558 1 2 404 320 4 2 19 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 160480 1 0 $X=20970 $Y=157520
X559 1 2 405 20 4 2 24 1 sky130_fd_sc_hd__dfrtp_4 $T=35880 171360 0 0 $X=35690 $Y=171120
X560 1 2 406 23 4 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=46920 149600 0 0 $X=46730 $Y=149360
X561 1 2 407 327 4 2 30 1 sky130_fd_sc_hd__dfrtp_4 $T=49220 171360 1 0 $X=49030 $Y=168400
X562 1 2 408 331 4 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=61640 160480 1 0 $X=61450 $Y=157520
X563 1 2 409 330 4 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=63020 160480 0 0 $X=62830 $Y=160240
X564 1 2 410 337 4 2 50 1 sky130_fd_sc_hd__dfrtp_4 $T=78660 160480 1 0 $X=78470 $Y=157520
X565 1 2 411 348 4 2 61 1 sky130_fd_sc_hd__dfrtp_4 $T=107640 160480 1 0 $X=107450 $Y=157520
X566 1 2 412 63 4 2 69 1 sky130_fd_sc_hd__dfrtp_4 $T=119140 149600 0 0 $X=118950 $Y=149360
X567 1 2 413 358 4 2 83 1 sky130_fd_sc_hd__dfrtp_4 $T=136160 160480 1 0 $X=135970 $Y=157520
X568 1 2 414 357 4 2 81 1 sky130_fd_sc_hd__dfrtp_4 $T=137080 155040 1 0 $X=136890 $Y=152080
X569 1 2 415 363 4 2 98 1 sky130_fd_sc_hd__dfrtp_4 $T=167440 171360 1 0 $X=167250 $Y=168400
X570 1 2 416 99 4 2 107 1 sky130_fd_sc_hd__dfrtp_4 $T=176180 171360 0 0 $X=175990 $Y=171120
X571 1 2 417 367 4 2 120 1 sky130_fd_sc_hd__dfrtp_4 $T=193200 171360 1 0 $X=193010 $Y=168400
X572 1 2 418 368 4 2 122 1 sky130_fd_sc_hd__dfrtp_4 $T=206080 165920 0 0 $X=205890 $Y=165680
X573 1 2 419 378 4 2 142 1 sky130_fd_sc_hd__dfrtp_4 $T=239660 155040 0 0 $X=239470 $Y=154800
X574 1 2 420 384 4 2 152 1 sky130_fd_sc_hd__dfrtp_4 $T=260360 149600 0 0 $X=260170 $Y=149360
X575 1 2 421 146 4 2 148 1 sky130_fd_sc_hd__dfrtp_4 $T=260820 171360 0 0 $X=260630 $Y=171120
X576 1 2 422 385 4 2 156 1 sky130_fd_sc_hd__dfrtp_4 $T=273700 160480 1 0 $X=273510 $Y=157520
X577 1 2 423 387 4 2 158 1 sky130_fd_sc_hd__dfrtp_4 $T=276920 171360 1 0 $X=276730 $Y=168400
X578 1 2 424 401 4 2 402 1 sky130_fd_sc_hd__dfrtp_4 $T=323840 160480 0 0 $X=323650 $Y=160240
X579 1 2 3 120 4 2 184 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 160480 1 0 $X=334690 $Y=157520
X580 1 2 3 402 4 2 185 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 165920 1 0 $X=334690 $Y=162960
X581 1 2 3 182 4 2 186 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 171360 1 0 $X=334690 $Y=168400
X582 1 2 22 ICV_13 $T=37260 160480 1 0 $X=37070 $Y=157520
X583 1 2 25 ICV_13 $T=45540 160480 0 0 $X=45350 $Y=160240
X584 1 2 340 ICV_13 $T=86020 160480 0 0 $X=85830 $Y=160240
X585 1 2 42 ICV_13 $T=90160 165920 0 0 $X=89970 $Y=165680
X586 1 2 353 ICV_13 $T=114080 155040 0 0 $X=113890 $Y=154800
X587 1 2 356 ICV_13 $T=132480 160480 1 0 $X=132290 $Y=157520
X588 1 2 76 ICV_13 $T=134780 165920 1 0 $X=134590 $Y=162960
X589 1 2 360 ICV_13 $T=154560 160480 1 0 $X=154370 $Y=157520
X590 1 2 90 ICV_13 $T=155480 165920 0 0 $X=155290 $Y=165680
X591 1 2 98 ICV_13 $T=170200 165920 0 0 $X=170010 $Y=165680
X592 1 2 110 ICV_13 $T=186760 171360 0 0 $X=186570 $Y=171120
X593 1 2 4 ICV_13 $T=202400 165920 0 0 $X=202210 $Y=165680
X594 1 2 118 ICV_13 $T=216660 165920 0 0 $X=216470 $Y=165680
X595 1 2 128 ICV_13 $T=235980 149600 0 0 $X=235790 $Y=149360
X596 1 2 380 ICV_13 $T=250240 165920 1 0 $X=250050 $Y=162960
X597 1 2 160 ICV_13 $T=282440 160480 0 0 $X=282250 $Y=160240
X598 1 2 389 ICV_13 $T=282440 165920 0 0 $X=282250 $Y=165680
X599 1 2 158 ICV_13 $T=282440 171360 0 0 $X=282250 $Y=171120
X600 1 2 164 ICV_13 $T=287500 171360 1 0 $X=287310 $Y=168400
X601 1 2 151 ICV_13 $T=294860 149600 0 0 $X=294670 $Y=149360
X602 1 2 166 ICV_13 $T=296240 165920 0 0 $X=296050 $Y=165680
X603 1 2 119 ICV_13 $T=301300 165920 0 0 $X=301110 $Y=165680
X604 1 2 110 ICV_13 $T=315100 165920 1 0 $X=314910 $Y=162960
X605 1 2 4 ICV_13 $T=320160 160480 0 0 $X=319970 $Y=160240
X606 1 2 170 ICV_13 $T=327520 149600 0 0 $X=327330 $Y=149360
X607 1 319 ICV_15 $T=17940 160480 1 0 $X=17750 $Y=157520
X608 1 19 ICV_15 $T=31740 155040 0 0 $X=31550 $Y=154800
X609 1 328 ICV_15 $T=46000 160480 1 0 $X=45810 $Y=157520
X610 1 328 ICV_15 $T=46000 165920 1 0 $X=45810 $Y=162960
X611 1 4 ICV_15 $T=59800 160480 0 0 $X=59610 $Y=160240
X612 1 50 ICV_15 $T=87860 155040 0 0 $X=87670 $Y=154800
X613 1 345 ICV_15 $T=102120 165920 1 0 $X=101930 $Y=162960
X614 1 346 ICV_15 $T=102120 171360 1 0 $X=101930 $Y=168400
X615 1 4 ICV_15 $T=115920 149600 0 0 $X=115730 $Y=149360
X616 1 67 ICV_15 $T=130180 165920 1 0 $X=129990 $Y=162960
X617 1 72 ICV_15 $T=130180 171360 1 0 $X=129990 $Y=168400
X618 1 81 ICV_15 $T=143980 149600 0 0 $X=143790 $Y=149360
X619 1 75 ICV_15 $T=143980 155040 0 0 $X=143790 $Y=154800
X620 1 82 ICV_15 $T=143980 171360 0 0 $X=143790 $Y=171120
X621 1 92 ICV_15 $T=158240 165920 1 0 $X=158050 $Y=162960
X622 1 91 ICV_15 $T=158240 171360 1 0 $X=158050 $Y=168400
X623 1 124 ICV_15 $T=214360 171360 1 0 $X=214170 $Y=168400
X624 1 136 ICV_15 $T=228160 160480 0 0 $X=227970 $Y=160240
X625 1 384 ICV_15 $T=256220 149600 0 0 $X=256030 $Y=149360
X626 1 48 ICV_15 $T=256220 160480 0 0 $X=256030 $Y=160240
X627 1 156 ICV_15 $T=284280 155040 0 0 $X=284090 $Y=154800
X628 1 168 ICV_15 $T=298540 155040 1 0 $X=298350 $Y=152080
X629 1 174 ICV_15 $T=312340 149600 0 0 $X=312150 $Y=149360
X630 1 2 318 ICV_16 $T=10120 165920 1 0 $X=9930 $Y=162960
X631 1 2 6 ICV_16 $T=11500 160480 1 0 $X=11310 $Y=157520
X632 1 2 325 ICV_16 $T=39100 165920 1 0 $X=38910 $Y=162960
X633 1 2 33 ICV_16 $T=68080 171360 1 0 $X=67890 $Y=168400
X634 1 2 352 ICV_16 $T=121440 155040 1 0 $X=121250 $Y=152080
X635 1 2 66 ICV_16 $T=121440 165920 0 0 $X=121250 $Y=165680
X636 1 2 61 ICV_16 $T=122820 160480 0 0 $X=122630 $Y=160240
X637 1 2 355 ICV_16 $T=152260 160480 0 0 $X=152070 $Y=160240
X638 1 2 13 ICV_16 $T=174340 155040 1 0 $X=174150 $Y=152080
X639 1 2 73 ICV_16 $T=181240 160480 0 0 $X=181050 $Y=160240
X640 1 2 84 ICV_16 $T=181700 155040 1 0 $X=181510 $Y=152080
X641 1 2 105 ICV_16 $T=181700 165920 0 0 $X=181510 $Y=165680
X642 1 2 121 ICV_16 $T=205620 155040 0 0 $X=205430 $Y=154800
X643 1 2 121 ICV_16 $T=205620 171360 0 0 $X=205430 $Y=171120
X644 1 2 67 ICV_16 $T=219420 149600 0 0 $X=219230 $Y=149360
X645 1 2 369 ICV_16 $T=220340 155040 0 0 $X=220150 $Y=154800
X646 1 2 142 ICV_16 $T=244720 149600 0 0 $X=244530 $Y=149360
X647 1 2 136 ICV_16 $T=251620 171360 0 0 $X=251430 $Y=171120
X648 1 2 148 ICV_16 $T=264500 165920 0 0 $X=264310 $Y=165680
X649 1 2 48 ICV_16 $T=265880 160480 0 0 $X=265690 $Y=160240
X650 1 2 392 ICV_16 $T=291180 155040 0 0 $X=290990 $Y=154800
X651 1 2 391 ICV_16 $T=292100 160480 1 0 $X=291910 $Y=157520
X652 1 2 160 ICV_16 $T=294860 160480 0 0 $X=294670 $Y=160240
X653 1 2 398 ICV_16 $T=316020 171360 1 0 $X=315830 $Y=168400
X654 1 2 399 ICV_16 $T=326140 155040 0 0 $X=325950 $Y=154800
X655 1 2 12 2 321 1 sky130_fd_sc_hd__inv_8 $T=21160 155040 0 0 $X=20970 $Y=154800
X656 1 2 19 2 325 1 sky130_fd_sc_hd__inv_8 $T=34960 155040 0 0 $X=34770 $Y=154800
X657 1 2 30 2 328 1 sky130_fd_sc_hd__inv_8 $T=53820 171360 0 0 $X=53630 $Y=171120
X658 1 2 36 2 334 1 sky130_fd_sc_hd__inv_8 $T=68080 165920 1 0 $X=67890 $Y=162960
X659 1 2 37 2 335 1 sky130_fd_sc_hd__inv_8 $T=71760 155040 0 0 $X=71570 $Y=154800
X660 1 2 50 2 340 1 sky130_fd_sc_hd__inv_8 $T=91080 155040 0 0 $X=90890 $Y=154800
X661 1 2 57 2 343 1 sky130_fd_sc_hd__inv_8 $T=103500 149600 0 0 $X=103310 $Y=149360
X662 1 2 61 2 345 1 sky130_fd_sc_hd__inv_8 $T=109940 160480 0 0 $X=109750 $Y=160240
X663 1 2 81 2 360 1 sky130_fd_sc_hd__inv_8 $T=147200 149600 0 0 $X=147010 $Y=149360
X664 1 2 83 2 355 1 sky130_fd_sc_hd__inv_8 $T=150420 160480 1 0 $X=150230 $Y=157520
X665 1 2 98 2 365 1 sky130_fd_sc_hd__inv_8 $T=175260 165920 0 0 $X=175070 $Y=165680
X666 1 2 122 2 369 1 sky130_fd_sc_hd__inv_8 $T=208380 165920 1 0 $X=208190 $Y=162960
X667 1 2 134 2 135 1 sky130_fd_sc_hd__inv_8 $T=225860 155040 1 0 $X=225670 $Y=152080
X668 1 2 142 2 375 1 sky130_fd_sc_hd__inv_8 $T=245640 155040 1 0 $X=245450 $Y=152080
X669 1 2 148 2 380 1 sky130_fd_sc_hd__inv_8 $T=264500 171360 1 0 $X=264310 $Y=168400
X670 1 2 156 2 389 1 sky130_fd_sc_hd__inv_8 $T=287040 160480 1 0 $X=286850 $Y=157520
X671 1 2 158 2 391 1 sky130_fd_sc_hd__inv_8 $T=287500 171360 0 0 $X=287310 $Y=171120
X672 1 2 173 2 394 1 sky130_fd_sc_hd__inv_8 $T=306360 171360 0 0 $X=306170 $Y=171120
X673 1 2 402 2 400 1 sky130_fd_sc_hd__inv_8 $T=327980 165920 0 0 $X=327790 $Y=165680
X674 1 2 11 319 2 318 1 sky130_fd_sc_hd__nor2_4 $T=21160 165920 1 0 $X=20970 $Y=162960
X675 1 2 16 322 2 320 1 sky130_fd_sc_hd__nor2_4 $T=25760 160480 0 0 $X=25570 $Y=160240
X676 1 2 16 326 2 327 1 sky130_fd_sc_hd__nor2_4 $T=40020 171360 1 0 $X=39830 $Y=168400
X677 1 2 33 332 2 330 1 sky130_fd_sc_hd__nor2_4 $T=66240 165920 0 0 $X=66050 $Y=165680
X678 1 2 33 333 2 331 1 sky130_fd_sc_hd__nor2_4 $T=68080 155040 1 0 $X=67890 $Y=152080
X679 1 2 338 336 2 337 1 sky130_fd_sc_hd__nor2_4 $T=81880 160480 0 0 $X=81690 $Y=160240
X680 1 2 338 342 2 56 1 sky130_fd_sc_hd__nor2_4 $T=95680 155040 1 0 $X=95490 $Y=152080
X681 1 2 338 58 2 59 1 sky130_fd_sc_hd__nor2_4 $T=104420 171360 0 0 $X=104230 $Y=171120
X682 1 2 338 346 2 348 1 sky130_fd_sc_hd__nor2_4 $T=105340 171360 1 0 $X=105150 $Y=168400
X683 1 2 338 350 2 63 1 sky130_fd_sc_hd__nor2_4 $T=109940 155040 0 0 $X=109750 $Y=154800
X684 1 2 70 354 2 358 1 sky130_fd_sc_hd__nor2_4 $T=136620 165920 0 0 $X=136430 $Y=165680
X685 1 2 70 356 2 357 1 sky130_fd_sc_hd__nor2_4 $T=138000 160480 0 0 $X=137810 $Y=160240
X686 1 2 70 362 2 363 1 sky130_fd_sc_hd__nor2_4 $T=151340 165920 0 0 $X=151150 $Y=165680
X687 1 2 106 113 2 367 1 sky130_fd_sc_hd__nor2_4 $T=190440 171360 0 0 $X=190250 $Y=171120
X688 1 2 106 114 2 115 1 sky130_fd_sc_hd__nor2_4 $T=191360 149600 0 0 $X=191170 $Y=149360
X689 1 2 125 371 2 126 1 sky130_fd_sc_hd__nor2_4 $T=216200 171360 0 0 $X=216010 $Y=171120
X690 1 2 125 370 2 368 1 sky130_fd_sc_hd__nor2_4 $T=217580 165920 1 0 $X=217390 $Y=162960
X691 1 2 139 376 2 378 1 sky130_fd_sc_hd__nor2_4 $T=235520 160480 1 0 $X=235330 $Y=157520
X692 1 2 125 383 2 146 1 sky130_fd_sc_hd__nor2_4 $T=254380 171360 1 0 $X=254190 $Y=168400
X693 1 2 125 382 2 384 1 sky130_fd_sc_hd__nor2_4 $T=259440 155040 0 0 $X=259250 $Y=154800
X694 1 2 154 386 2 385 1 sky130_fd_sc_hd__nor2_4 $T=278300 160480 0 0 $X=278110 $Y=160240
X695 1 2 154 388 2 387 1 sky130_fd_sc_hd__nor2_4 $T=278300 165920 0 0 $X=278110 $Y=165680
X696 1 2 170 395 2 177 1 sky130_fd_sc_hd__nor2_4 $T=306360 155040 0 0 $X=306170 $Y=154800
X697 1 2 170 397 2 172 1 sky130_fd_sc_hd__nor2_4 $T=308660 171360 1 0 $X=308470 $Y=168400
X698 1 2 170 398 2 401 1 sky130_fd_sc_hd__nor2_4 $T=316020 160480 0 0 $X=315830 $Y=160240
X699 1 2 170 180 2 181 1 sky130_fd_sc_hd__nor2_4 $T=331200 149600 0 0 $X=331010 $Y=149360
X700 1 2 321 7 10 323 2 319 1 sky130_fd_sc_hd__o22a_4 $T=23000 171360 1 0 $X=22810 $Y=168400
X701 1 2 325 22 21 324 2 322 1 sky130_fd_sc_hd__o22a_4 $T=39100 160480 0 0 $X=38910 $Y=160240
X702 1 2 328 22 21 329 2 326 1 sky130_fd_sc_hd__o22a_4 $T=49220 165920 1 0 $X=49030 $Y=162960
X703 1 2 334 38 39 45 2 332 1 sky130_fd_sc_hd__o22a_4 $T=74520 171360 0 0 $X=74330 $Y=171120
X704 1 2 335 43 41 339 2 333 1 sky130_fd_sc_hd__o22a_4 $T=79120 149600 0 0 $X=78930 $Y=149360
X705 1 2 340 51 52 341 2 336 1 sky130_fd_sc_hd__o22a_4 $T=90620 165920 1 0 $X=90430 $Y=162960
X706 1 2 343 51 52 344 2 342 1 sky130_fd_sc_hd__o22a_4 $T=95680 160480 0 0 $X=95490 $Y=160240
X707 1 2 345 51 52 347 2 346 1 sky130_fd_sc_hd__o22a_4 $T=105340 165920 1 0 $X=105150 $Y=162960
X708 1 2 62 351 353 349 2 58 1 sky130_fd_sc_hd__o22a_4 $T=112240 171360 1 0 $X=112050 $Y=168400
X709 1 2 60 351 353 352 2 350 1 sky130_fd_sc_hd__o22a_4 $T=119140 155040 0 0 $X=118950 $Y=154800
X710 1 2 355 29 31 359 2 354 1 sky130_fd_sc_hd__o22a_4 $T=138460 165920 1 0 $X=138270 $Y=162960
X711 1 2 360 80 75 361 2 356 1 sky130_fd_sc_hd__o22a_4 $T=147200 155040 0 0 $X=147010 $Y=154800
X712 1 2 91 92 90 364 2 93 1 sky130_fd_sc_hd__o22a_4 $T=159160 165920 0 0 $X=158970 $Y=165680
X713 1 2 365 92 90 366 2 362 1 sky130_fd_sc_hd__o22a_4 $T=164680 165920 1 0 $X=164490 $Y=162960
X714 1 2 369 351 353 372 2 370 1 sky130_fd_sc_hd__o22a_4 $T=211600 160480 0 0 $X=211410 $Y=160240
X715 1 2 129 130 131 373 2 371 1 sky130_fd_sc_hd__o22a_4 $T=222180 171360 1 0 $X=221990 $Y=168400
X716 1 2 375 130 131 374 2 376 1 sky130_fd_sc_hd__o22a_4 $T=234140 165920 1 0 $X=233950 $Y=162960
X717 1 2 141 130 131 377 2 140 1 sky130_fd_sc_hd__o22a_4 $T=240580 171360 0 0 $X=240390 $Y=171120
X718 1 2 144 351 353 381 2 382 1 sky130_fd_sc_hd__o22a_4 $T=253000 160480 1 0 $X=252810 $Y=157520
X719 1 2 380 351 353 379 2 383 1 sky130_fd_sc_hd__o22a_4 $T=253920 165920 1 0 $X=253730 $Y=162960
X720 1 2 391 157 160 392 2 388 1 sky130_fd_sc_hd__o22a_4 $T=287040 165920 1 0 $X=286850 $Y=162960
X721 1 2 389 157 160 390 2 386 1 sky130_fd_sc_hd__o22a_4 $T=287500 160480 0 0 $X=287310 $Y=160240
X722 1 2 394 174 176 393 2 397 1 sky130_fd_sc_hd__o22a_4 $T=308660 165920 1 0 $X=308470 $Y=162960
X723 1 2 175 174 176 396 2 395 1 sky130_fd_sc_hd__o22a_4 $T=310500 155040 1 0 $X=310310 $Y=152080
X724 1 2 400 174 176 399 2 398 1 sky130_fd_sc_hd__o22a_4 $T=318320 160480 1 0 $X=318130 $Y=157520
X725 1 2 178 174 176 179 2 180 1 sky130_fd_sc_hd__o22a_4 $T=321080 149600 0 0 $X=320890 $Y=149360
X726 1 2 29 2 22 1 sky130_fd_sc_hd__buf_1 $T=53820 155040 0 0 $X=53630 $Y=154800
X727 1 2 31 2 21 1 sky130_fd_sc_hd__buf_1 $T=56120 160480 1 0 $X=55930 $Y=157520
X728 1 2 35 2 33 1 sky130_fd_sc_hd__buf_1 $T=66700 171360 0 0 $X=66510 $Y=171120
X729 1 2 44 2 11 1 sky130_fd_sc_hd__buf_1 $T=79580 171360 1 0 $X=79390 $Y=168400
X730 1 2 44 2 338 1 sky130_fd_sc_hd__buf_1 $T=96600 171360 0 0 $X=96410 $Y=171120
X731 1 2 55 2 40 1 sky130_fd_sc_hd__buf_1 $T=97520 171360 1 0 $X=97330 $Y=168400
X732 1 2 66 2 53 1 sky130_fd_sc_hd__buf_1 $T=119140 165920 0 0 $X=118950 $Y=165680
X733 1 2 67 2 35 1 sky130_fd_sc_hd__buf_1 $T=126500 171360 0 0 $X=126310 $Y=171120
X734 1 2 55 2 71 1 sky130_fd_sc_hd__buf_1 $T=131560 165920 0 0 $X=131370 $Y=165680
X735 1 2 55 2 13 1 sky130_fd_sc_hd__buf_1 $T=133400 165920 1 0 $X=133210 $Y=162960
X736 1 2 67 2 44 1 sky130_fd_sc_hd__buf_1 $T=133400 171360 1 0 $X=133210 $Y=168400
X737 1 2 77 2 29 1 sky130_fd_sc_hd__buf_1 $T=137540 149600 0 0 $X=137350 $Y=149360
X738 1 2 74 2 31 1 sky130_fd_sc_hd__buf_1 $T=140300 155040 0 0 $X=140110 $Y=154800
X739 1 2 67 2 84 1 sky130_fd_sc_hd__buf_1 $T=147200 165920 0 0 $X=147010 $Y=165680
X740 1 2 55 2 88 1 sky130_fd_sc_hd__buf_1 $T=161460 171360 1 0 $X=161270 $Y=168400
X741 1 2 87 2 101 1 sky130_fd_sc_hd__buf_1 $T=174800 165920 1 0 $X=174610 $Y=162960
X742 1 2 102 2 55 1 sky130_fd_sc_hd__buf_1 $T=176640 160480 1 0 $X=176450 $Y=157520
X743 1 2 73 2 103 1 sky130_fd_sc_hd__buf_1 $T=178940 160480 0 0 $X=178750 $Y=160240
X744 1 2 89 2 104 1 sky130_fd_sc_hd__buf_1 $T=180320 155040 0 0 $X=180130 $Y=154800
X745 1 2 84 2 106 1 sky130_fd_sc_hd__buf_1 $T=181700 160480 1 0 $X=181510 $Y=157520
X746 1 2 105 2 92 1 sky130_fd_sc_hd__buf_1 $T=181700 171360 1 0 $X=181510 $Y=168400
X747 1 2 108 2 109 1 sky130_fd_sc_hd__buf_1 $T=185380 155040 0 0 $X=185190 $Y=154800
X748 1 2 102 2 66 1 sky130_fd_sc_hd__buf_1 $T=190440 160480 1 0 $X=190250 $Y=157520
X749 1 2 111 2 112 1 sky130_fd_sc_hd__buf_1 $T=191360 155040 0 0 $X=191170 $Y=154800
X750 1 2 79 2 110 1 sky130_fd_sc_hd__buf_1 $T=192280 165920 0 0 $X=192090 $Y=165680
X751 1 2 85 2 117 1 sky130_fd_sc_hd__buf_1 $T=196880 155040 0 0 $X=196690 $Y=154800
X752 1 2 118 2 119 1 sky130_fd_sc_hd__buf_1 $T=198720 165920 1 0 $X=198530 $Y=162960
X753 1 2 121 2 67 1 sky130_fd_sc_hd__buf_1 $T=205620 160480 1 0 $X=205430 $Y=157520
X754 1 2 66 2 123 1 sky130_fd_sc_hd__buf_1 $T=207460 171360 1 0 $X=207270 $Y=168400
X755 1 2 67 2 128 1 sky130_fd_sc_hd__buf_1 $T=217120 149600 0 0 $X=216930 $Y=149360
X756 1 2 132 2 105 1 sky130_fd_sc_hd__buf_1 $T=224480 165920 1 0 $X=224290 $Y=162960
X757 1 2 138 2 97 1 sky130_fd_sc_hd__buf_1 $T=232300 171360 1 0 $X=232110 $Y=168400
X758 1 2 132 2 130 1 sky130_fd_sc_hd__buf_1 $T=233220 165920 0 0 $X=233030 $Y=165680
X759 1 2 132 2 351 1 sky130_fd_sc_hd__buf_1 $T=233680 155040 0 0 $X=233490 $Y=154800
X760 1 2 128 2 125 1 sky130_fd_sc_hd__buf_1 $T=237820 155040 1 0 $X=237630 $Y=152080
X761 1 2 138 2 131 1 sky130_fd_sc_hd__buf_1 $T=241040 165920 0 0 $X=240850 $Y=165680
X762 1 2 138 2 353 1 sky130_fd_sc_hd__buf_1 $T=248860 160480 0 0 $X=248670 $Y=160240
X763 1 2 65 2 147 1 sky130_fd_sc_hd__buf_1 $T=259440 165920 0 0 $X=259250 $Y=165680
X764 1 2 64 2 149 1 sky130_fd_sc_hd__buf_1 $T=265420 155040 1 0 $X=265230 $Y=152080
X765 1 2 48 2 150 1 sky130_fd_sc_hd__buf_1 $T=265880 165920 1 0 $X=265690 $Y=162960
X766 1 2 127 2 151 1 sky130_fd_sc_hd__buf_1 $T=266340 155040 0 0 $X=266150 $Y=154800
X767 1 2 145 2 153 1 sky130_fd_sc_hd__buf_1 $T=274620 149600 0 0 $X=274430 $Y=149360
X768 1 2 166 2 159 1 sky130_fd_sc_hd__buf_1 $T=299920 165920 0 0 $X=299730 $Y=165680
X769 1 2 169 2 160 1 sky130_fd_sc_hd__buf_1 $T=301760 155040 1 0 $X=301570 $Y=152080
X770 1 2 166 2 171 1 sky130_fd_sc_hd__buf_1 $T=303600 165920 1 0 $X=303410 $Y=162960
X771 1 2 15 17 13 2 14 1 sky130_fd_sc_hd__o21a_4 $T=24380 171360 0 0 $X=24190 $Y=171120
X772 1 2 18 321 13 2 323 1 sky130_fd_sc_hd__o21a_4 $T=28060 165920 1 0 $X=27870 $Y=162960
X773 1 2 26 328 27 2 329 1 sky130_fd_sc_hd__o21a_4 $T=47380 165920 0 0 $X=47190 $Y=165680
X774 1 2 25 325 27 2 324 1 sky130_fd_sc_hd__o21a_4 $T=49220 160480 0 0 $X=49030 $Y=160240
X775 1 2 42 334 40 2 45 1 sky130_fd_sc_hd__o21a_4 $T=80040 165920 0 0 $X=79850 $Y=165680
X776 1 2 48 335 40 2 339 1 sky130_fd_sc_hd__o21a_4 $T=84180 155040 1 0 $X=83990 $Y=152080
X777 1 2 49 46 40 2 47 1 sky130_fd_sc_hd__o21a_4 $T=84640 171360 1 0 $X=84450 $Y=168400
X778 1 2 42 340 53 2 341 1 sky130_fd_sc_hd__o21a_4 $T=93840 165920 0 0 $X=93650 $Y=165680
X779 1 2 54 343 53 2 344 1 sky130_fd_sc_hd__o21a_4 $T=98440 155040 0 0 $X=98250 $Y=154800
X780 1 2 49 345 53 2 347 1 sky130_fd_sc_hd__o21a_4 $T=105340 165920 0 0 $X=105150 $Y=165680
X781 1 2 65 62 53 2 349 1 sky130_fd_sc_hd__o21a_4 $T=114540 165920 1 0 $X=114350 $Y=162960
X782 1 2 64 60 53 2 352 1 sky130_fd_sc_hd__o21a_4 $T=115000 155040 1 0 $X=114810 $Y=152080
X783 1 2 73 72 71 2 68 1 sky130_fd_sc_hd__o21a_4 $T=133400 171360 0 0 $X=133210 $Y=171120
X784 1 2 79 76 71 2 78 1 sky130_fd_sc_hd__o21a_4 $T=137540 171360 1 0 $X=137350 $Y=168400
X785 1 2 85 355 88 2 359 1 sky130_fd_sc_hd__o21a_4 $T=148580 165920 1 0 $X=148390 $Y=162960
X786 1 2 87 82 88 2 86 1 sky130_fd_sc_hd__o21a_4 $T=151800 171360 0 0 $X=151610 $Y=171120
X787 1 2 89 360 88 2 361 1 sky130_fd_sc_hd__o21a_4 $T=156400 155040 0 0 $X=156210 $Y=154800
X788 1 2 94 91 88 2 364 1 sky130_fd_sc_hd__o21a_4 $T=161920 171360 0 0 $X=161730 $Y=171120
X789 1 2 95 365 88 2 366 1 sky130_fd_sc_hd__o21a_4 $T=164680 160480 0 0 $X=164490 $Y=160240
X790 1 2 25 96 13 2 100 1 sky130_fd_sc_hd__o21a_4 $T=175260 149600 0 0 $X=175070 $Y=149360
X791 1 2 127 369 123 2 372 1 sky130_fd_sc_hd__o21a_4 $T=217580 160480 1 0 $X=217390 $Y=157520
X792 1 2 118 129 123 2 373 1 sky130_fd_sc_hd__o21a_4 $T=220340 165920 0 0 $X=220150 $Y=165680
X793 1 2 89 375 136 2 374 1 sky130_fd_sc_hd__o21a_4 $T=231840 160480 0 0 $X=231650 $Y=160240
X794 1 2 79 141 123 2 377 1 sky130_fd_sc_hd__o21a_4 $T=245640 171360 1 0 $X=245450 $Y=168400
X795 1 2 145 144 123 2 381 1 sky130_fd_sc_hd__o21a_4 $T=256220 155040 1 0 $X=256030 $Y=152080
X796 1 2 48 380 123 2 379 1 sky130_fd_sc_hd__o21a_4 $T=259440 160480 0 0 $X=259250 $Y=160240
X797 1 2 149 162 159 2 161 1 sky130_fd_sc_hd__o21a_4 $T=289340 149600 0 0 $X=289150 $Y=149360
X798 1 2 153 155 159 2 163 1 sky130_fd_sc_hd__o21a_4 $T=289340 155040 1 0 $X=289150 $Y=152080
X799 1 2 150 391 159 2 392 1 sky130_fd_sc_hd__o21a_4 $T=290720 165920 0 0 $X=290530 $Y=165680
X800 1 2 147 389 164 2 390 1 sky130_fd_sc_hd__o21a_4 $T=291180 171360 1 0 $X=290990 $Y=168400
X801 1 2 151 168 159 2 167 1 sky130_fd_sc_hd__o21a_4 $T=298540 149600 0 0 $X=298350 $Y=149360
X802 1 2 119 394 159 2 393 1 sky130_fd_sc_hd__o21a_4 $T=304980 165920 0 0 $X=304790 $Y=165680
X803 1 2 101 175 171 2 396 1 sky130_fd_sc_hd__o21a_4 $T=309120 160480 1 0 $X=308930 $Y=157520
X804 1 2 110 400 171 2 399 1 sky130_fd_sc_hd__o21a_4 $T=318780 165920 1 0 $X=318590 $Y=162960
X805 1 2 103 178 171 2 179 1 sky130_fd_sc_hd__o21a_4 $T=319700 155040 0 0 $X=319510 $Y=154800
X806 1 2 ICV_23 $T=6900 149600 0 0 $X=6710 $Y=149360
X807 1 2 ICV_23 $T=6900 171360 1 0 $X=6710 $Y=168400
X808 1 2 ICV_23 $T=17940 149600 0 0 $X=17750 $Y=149360
X809 1 2 ICV_23 $T=23920 155040 1 0 $X=23730 $Y=152080
X810 1 2 ICV_23 $T=34960 155040 1 0 $X=34770 $Y=152080
X811 1 2 ICV_23 $T=48300 155040 1 0 $X=48110 $Y=152080
X812 1 2 ICV_23 $T=151340 149600 0 0 $X=151150 $Y=149360
X813 1 2 ICV_23 $T=160540 155040 1 0 $X=160350 $Y=152080
X814 1 2 ICV_23 $T=161920 155040 0 0 $X=161730 $Y=154800
X815 1 2 ICV_23 $T=176180 165920 1 0 $X=175990 $Y=162960
X816 1 2 ICV_23 $T=187680 160480 0 0 $X=187490 $Y=160240
X817 1 2 ICV_23 $T=188600 155040 1 0 $X=188410 $Y=152080
X818 1 2 ICV_23 $T=191820 160480 1 0 $X=191630 $Y=157520
X819 1 2 ICV_23 $T=199640 155040 1 0 $X=199450 $Y=152080
X820 1 2 ICV_23 $T=202400 149600 0 0 $X=202210 $Y=149360
X821 1 2 ICV_23 $T=271400 171360 0 0 $X=271210 $Y=171120
X822 1 2 ICV_23 $T=272780 155040 1 0 $X=272590 $Y=152080
X823 1 2 ICV_23 $T=314640 171360 0 0 $X=314450 $Y=171120
X824 1 2 ICV_23 $T=328900 155040 1 0 $X=328710 $Y=152080
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or2_4 VNB VPB B A VPWR X VGND
** N=37 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 8 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1740 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2580 $Y=235 $D=9
M6 9 B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=455 $Y=1485 $D=89
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2160 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176
** N=422 EP=176 IP=3559 FDC=4555
*.SEEDPROM
X0 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=129145 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=134585 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=140025 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=145465 $D=191
X4 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 127840 1 0 $X=5330 $Y=124880
X5 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 127840 0 0 $X=5330 $Y=127600
X6 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 133280 1 0 $X=5330 $Y=130320
X7 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 133280 0 0 $X=5330 $Y=133040
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 138720 1 0 $X=5330 $Y=135760
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 138720 0 0 $X=5330 $Y=138480
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 144160 1 0 $X=5330 $Y=141200
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 144160 0 0 $X=5330 $Y=143920
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 149600 1 0 $X=5330 $Y=146640
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 127840 1 0 $X=6710 $Y=124880
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 127840 0 0 $X=6710 $Y=127600
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 133280 1 0 $X=6710 $Y=130320
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 127840 1 0 $X=18210 $Y=124880
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=23920 127840 1 0 $X=23730 $Y=124880
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 133280 1 0 $X=25570 $Y=130320
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28520 127840 0 0 $X=28330 $Y=127600
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=46460 133280 1 0 $X=46270 $Y=130320
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=67160 149600 1 0 $X=66970 $Y=146640
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 144160 1 0 $X=76170 $Y=141200
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=83260 149600 1 0 $X=83070 $Y=146640
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88320 133280 0 0 $X=88130 $Y=133040
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88780 138720 1 0 $X=88590 $Y=135760
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 144160 1 0 $X=102390 $Y=141200
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=113620 149600 1 0 $X=113430 $Y=146640
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=141680 149600 1 0 $X=141490 $Y=146640
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 127840 0 0 $X=144250 $Y=127600
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 127840 1 0 $X=158510 $Y=124880
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 149600 1 0 $X=158510 $Y=146640
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=168820 144160 0 0 $X=168630 $Y=143920
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=172500 127840 0 0 $X=172310 $Y=127600
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=186760 133280 1 0 $X=186570 $Y=130320
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=194580 144160 0 0 $X=194390 $Y=143920
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 144160 1 0 $X=214630 $Y=141200
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224940 133280 0 0 $X=224750 $Y=133040
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=238280 127840 1 0 $X=238090 $Y=124880
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=250240 133280 1 0 $X=250050 $Y=130320
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=250240 133280 0 0 $X=250050 $Y=133040
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=251620 138720 0 0 $X=251430 $Y=138480
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=256220 127840 1 0 $X=256030 $Y=124880
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=257140 133280 1 0 $X=256950 $Y=130320
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 133280 1 0 $X=270750 $Y=130320
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=302220 133280 0 0 $X=302030 $Y=133040
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=312800 127840 0 0 $X=312610 $Y=127600
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 133280 0 0 $X=314450 $Y=133040
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=315560 127840 1 0 $X=315370 $Y=124880
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=319700 127840 1 0 $X=319510 $Y=124880
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 138720 0 0 $X=340670 $Y=138480
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 144160 0 0 $X=340670 $Y=143920
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 127840 0 180 $X=348950 $Y=124880
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 127840 1 180 $X=348950 $Y=127600
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 133280 0 180 $X=348950 $Y=130320
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 133280 1 180 $X=348950 $Y=133040
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 138720 0 180 $X=348950 $Y=135760
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 138720 1 180 $X=348950 $Y=138480
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 144160 0 180 $X=348950 $Y=141200
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 144160 1 180 $X=348950 $Y=143920
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 149600 0 180 $X=348950 $Y=146640
X152 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=14720 127840 1 0 $X=14530 $Y=124880
X153 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 127840 1 0 $X=20050 $Y=124880
X154 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=33580 149600 1 0 $X=33390 $Y=146640
X155 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34960 144160 1 0 $X=34770 $Y=141200
X156 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 149600 1 0 $X=43970 $Y=146640
X157 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57040 127840 0 0 $X=56850 $Y=127600
X158 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=59340 138720 1 0 $X=59150 $Y=135760
X159 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=62100 144160 0 0 $X=61910 $Y=143920
X160 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71300 133280 1 0 $X=71110 $Y=130320
X161 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71760 138720 1 0 $X=71570 $Y=135760
X162 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 127840 1 0 $X=72030 $Y=124880
X163 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 138720 1 0 $X=76170 $Y=135760
X164 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=85100 138720 1 0 $X=84910 $Y=135760
X165 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=98900 144160 1 0 $X=98710 $Y=141200
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=115460 144160 1 0 $X=115270 $Y=141200
X167 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 138720 1 0 $X=128150 $Y=135760
X168 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=130640 138720 0 0 $X=130450 $Y=138480
X169 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 138720 1 0 $X=132290 $Y=135760
X170 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 144160 1 0 $X=132290 $Y=141200
X171 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 133280 1 0 $X=139650 $Y=130320
X172 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=155020 127840 1 0 $X=154830 $Y=124880
X173 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=157320 133280 0 0 $X=157130 $Y=133040
X174 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=162380 127840 1 0 $X=162190 $Y=124880
X175 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165140 149600 1 0 $X=164950 $Y=146640
X176 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 138720 1 0 $X=184270 $Y=135760
X177 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=187680 133280 0 0 $X=187490 $Y=133040
X178 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 127840 1 0 $X=188410 $Y=124880
X179 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 144160 1 0 $X=188410 $Y=141200
X180 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=192280 149600 1 0 $X=192090 $Y=146640
X181 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=192740 133280 0 0 $X=192550 $Y=133040
X182 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=196420 127840 0 0 $X=196230 $Y=127600
X183 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=197800 133280 0 0 $X=197610 $Y=133040
X184 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=209760 127840 1 0 $X=209570 $Y=124880
X185 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=223100 144160 0 0 $X=222910 $Y=143920
X186 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 133280 1 0 $X=240390 $Y=130320
X187 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=251620 138720 1 0 $X=251430 $Y=135760
X188 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=252540 127840 1 0 $X=252350 $Y=124880
X189 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=265420 127840 1 0 $X=265230 $Y=124880
X190 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267260 133280 1 0 $X=267070 $Y=130320
X191 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 149600 1 0 $X=268450 $Y=146640
X192 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 138720 1 0 $X=272590 $Y=135760
X193 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 138720 0 0 $X=272590 $Y=138480
X194 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 144160 1 0 $X=272590 $Y=141200
X195 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=279220 133280 0 0 $X=279030 $Y=133040
X196 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=309580 133280 0 0 $X=309390 $Y=133040
X197 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310960 144160 1 0 $X=310770 $Y=141200
X198 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=311880 127840 1 0 $X=311690 $Y=124880
X199 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=311880 138720 1 0 $X=311690 $Y=135760
X200 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314180 133280 1 0 $X=313990 $Y=130320
X201 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=323840 149600 1 0 $X=323650 $Y=146640
X202 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324300 144160 1 0 $X=324110 $Y=141200
X203 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=325220 138720 0 0 $X=325030 $Y=138480
X204 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 127840 1 0 $X=344810 $Y=124880
X205 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 138720 1 0 $X=344810 $Y=135760
X206 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 133280 1 0 $X=345270 $Y=130320
X207 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 149600 1 0 $X=345270 $Y=146640
X208 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=14260 149600 1 0 $X=14070 $Y=146640
X209 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=20240 133280 1 0 $X=20050 $Y=130320
X210 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40940 133280 1 0 $X=40750 $Y=130320
X211 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=48300 127840 1 0 $X=48110 $Y=124880
X212 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55660 144160 1 0 $X=55470 $Y=141200
X213 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=60260 127840 1 0 $X=60070 $Y=124880
X214 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=64860 133280 1 0 $X=64670 $Y=130320
X215 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=65780 138720 0 0 $X=65590 $Y=138480
X216 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=87400 133280 1 0 $X=87210 $Y=130320
X217 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=96600 138720 1 0 $X=96410 $Y=135760
X218 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=109480 127840 1 0 $X=109290 $Y=124880
X219 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=133860 144160 0 0 $X=133670 $Y=143920
X220 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=151340 144160 1 0 $X=151150 $Y=141200
X221 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=152260 138720 0 0 $X=152070 $Y=138480
X222 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=152720 144160 0 0 $X=152530 $Y=143920
X223 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=153640 138720 1 0 $X=153450 $Y=135760
X224 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=154100 133280 1 0 $X=153910 $Y=130320
X225 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=166980 127840 0 0 $X=166790 $Y=127600
X226 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=167440 127840 1 0 $X=167250 $Y=124880
X227 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=189060 144160 0 0 $X=188870 $Y=143920
X228 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=207460 127840 0 0 $X=207270 $Y=127600
X229 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=208840 133280 1 0 $X=208650 $Y=130320
X230 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=209300 144160 1 0 $X=209110 $Y=141200
X231 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=236900 149600 1 0 $X=236710 $Y=146640
X232 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=243800 127840 0 0 $X=243610 $Y=127600
X233 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=244720 133280 1 0 $X=244530 $Y=130320
X234 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=244720 144160 1 0 $X=244530 $Y=141200
X235 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=246100 138720 0 0 $X=245910 $Y=138480
X236 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=263580 144160 1 0 $X=263390 $Y=141200
X237 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=265880 138720 1 0 $X=265690 $Y=135760
X238 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=279220 127840 1 0 $X=279030 $Y=124880
X239 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=283820 133280 1 0 $X=283630 $Y=130320
X240 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293940 127840 1 0 $X=293750 $Y=124880
X241 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=294400 138720 1 0 $X=294210 $Y=135760
X242 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=302220 127840 0 0 $X=302030 $Y=127600
X243 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=318780 133280 0 0 $X=318590 $Y=133040
X244 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322920 133280 1 0 $X=322730 $Y=130320
X245 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=328900 127840 1 0 $X=328710 $Y=124880
X246 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=328900 133280 1 0 $X=328710 $Y=130320
X247 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=328900 138720 1 0 $X=328710 $Y=135760
X248 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=340400 144160 1 0 $X=340210 $Y=141200
X249 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=342700 127840 0 0 $X=342510 $Y=127600
X250 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=342700 133280 0 0 $X=342510 $Y=133040
X251 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=342700 138720 0 0 $X=342510 $Y=138480
X252 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=342700 144160 0 0 $X=342510 $Y=143920
X253 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=14260 133280 0 0 $X=14070 $Y=133040
X254 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18860 127840 0 0 $X=18670 $Y=127600
X255 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=22080 133280 0 0 $X=21890 $Y=133040
X256 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=25760 144160 0 0 $X=25570 $Y=143920
X257 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 144160 1 0 $X=31550 $Y=141200
X258 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=32200 127840 1 0 $X=32010 $Y=124880
X259 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=43700 138720 1 0 $X=43510 $Y=135760
X260 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=48300 133280 1 0 $X=48110 $Y=130320
X261 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=48300 138720 1 0 $X=48110 $Y=135760
X262 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=57960 133280 0 0 $X=57770 $Y=133040
X263 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=72220 144160 1 0 $X=72030 $Y=141200
X264 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=72680 144160 0 0 $X=72490 $Y=143920
X265 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=77280 138720 0 0 $X=77090 $Y=138480
X266 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=92920 133280 1 0 $X=92730 $Y=130320
X267 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 138720 1 0 $X=101930 $Y=135760
X268 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=105800 127840 0 0 $X=105610 $Y=127600
X269 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=105800 133280 0 0 $X=105610 $Y=133040
X270 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=113620 127840 0 0 $X=113430 $Y=127600
X271 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=113620 133280 0 0 $X=113430 $Y=133040
X272 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 138720 0 0 $X=118030 $Y=138480
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=126040 149600 1 0 $X=125850 $Y=146640
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=144440 149600 1 0 $X=144250 $Y=146640
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 133280 1 0 $X=160350 $Y=130320
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 149600 1 0 $X=160350 $Y=146640
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=162380 127840 0 0 $X=162190 $Y=127600
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=170200 138720 0 0 $X=170010 $Y=138480
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174800 133280 1 0 $X=174610 $Y=130320
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188140 138720 0 0 $X=187950 $Y=138480
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=193200 138720 1 0 $X=193010 $Y=135760
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=204700 144160 0 0 $X=204510 $Y=143920
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=206540 149600 1 0 $X=206350 $Y=146640
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=212980 127840 0 0 $X=212790 $Y=127600
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 133280 1 0 $X=214170 $Y=130320
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=215740 138720 0 0 $X=215550 $Y=138480
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 127840 1 0 $X=216470 $Y=124880
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 149600 1 0 $X=216470 $Y=146640
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=224940 138720 0 0 $X=224750 $Y=138480
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=225400 127840 1 0 $X=225210 $Y=124880
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226320 133280 1 0 $X=226130 $Y=130320
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230460 133280 0 0 $X=230270 $Y=133040
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=233220 144160 1 0 $X=233030 $Y=141200
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=235520 127840 1 0 $X=235330 $Y=124880
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=241960 144160 1 0 $X=241770 $Y=141200
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 149600 1 0 $X=242230 $Y=146640
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 144160 0 0 $X=258330 $Y=143920
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=281980 149600 1 0 $X=281790 $Y=146640
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=282440 144160 0 0 $X=282250 $Y=143920
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284740 127840 1 0 $X=284550 $Y=124880
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=289340 133280 1 0 $X=289150 $Y=130320
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298080 133280 1 0 $X=297890 $Y=130320
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=299920 138720 0 0 $X=299730 $Y=138480
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=303140 138720 1 0 $X=302950 $Y=135760
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=307740 127840 0 0 $X=307550 $Y=127600
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=318780 149600 1 0 $X=318590 $Y=146640
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 149600 1 0 $X=328710 $Y=146640
X308 1 312 sky130_fd_sc_hd__diode_2 $T=16100 133280 0 0 $X=15910 $Y=133040
X309 1 4 sky130_fd_sc_hd__diode_2 $T=19320 138720 0 0 $X=19130 $Y=138480
X310 1 7 sky130_fd_sc_hd__diode_2 $T=20700 127840 0 0 $X=20510 $Y=127600
X311 1 318 sky130_fd_sc_hd__diode_2 $T=26220 138720 1 0 $X=26030 $Y=135760
X312 1 315 sky130_fd_sc_hd__diode_2 $T=26220 138720 0 0 $X=26030 $Y=138480
X313 1 9 sky130_fd_sc_hd__diode_2 $T=27600 127840 0 0 $X=27410 $Y=127600
X314 1 320 sky130_fd_sc_hd__diode_2 $T=28980 127840 1 0 $X=28790 $Y=124880
X315 1 323 sky130_fd_sc_hd__diode_2 $T=34040 144160 1 0 $X=33850 $Y=141200
X316 1 325 sky130_fd_sc_hd__diode_2 $T=38180 149600 1 0 $X=37990 $Y=146640
X317 1 18 sky130_fd_sc_hd__diode_2 $T=41400 138720 0 0 $X=41210 $Y=138480
X318 1 29 sky130_fd_sc_hd__diode_2 $T=65320 127840 0 0 $X=65130 $Y=127600
X319 1 30 sky130_fd_sc_hd__diode_2 $T=66700 144160 0 0 $X=66510 $Y=143920
X320 1 334 sky130_fd_sc_hd__diode_2 $T=70380 133280 1 0 $X=70190 $Y=130320
X321 1 32 sky130_fd_sc_hd__diode_2 $T=71300 138720 0 0 $X=71110 $Y=138480
X322 1 336 sky130_fd_sc_hd__diode_2 $T=82340 149600 1 0 $X=82150 $Y=146640
X323 1 4 sky130_fd_sc_hd__diode_2 $T=93380 127840 0 0 $X=93190 $Y=127600
X324 1 4 sky130_fd_sc_hd__diode_2 $T=93380 133280 0 0 $X=93190 $Y=133040
X325 1 4 sky130_fd_sc_hd__diode_2 $T=96140 144160 0 0 $X=95950 $Y=143920
X326 1 46 sky130_fd_sc_hd__diode_2 $T=107640 127840 0 0 $X=107450 $Y=127600
X327 1 47 sky130_fd_sc_hd__diode_2 $T=107640 133280 0 0 $X=107450 $Y=133040
X328 1 53 sky130_fd_sc_hd__diode_2 $T=118220 149600 1 0 $X=118030 $Y=146640
X329 1 54 sky130_fd_sc_hd__diode_2 $T=119600 144160 1 0 $X=119410 $Y=141200
X330 1 59 sky130_fd_sc_hd__diode_2 $T=126500 144160 0 0 $X=126310 $Y=143920
X331 1 343 sky130_fd_sc_hd__diode_2 $T=127420 138720 1 0 $X=127230 $Y=135760
X332 1 342 sky130_fd_sc_hd__diode_2 $T=128340 149600 1 0 $X=128150 $Y=146640
X333 1 63 sky130_fd_sc_hd__diode_2 $T=130640 127840 0 0 $X=130450 $Y=127600
X334 1 345 sky130_fd_sc_hd__diode_2 $T=136160 138720 1 0 $X=135970 $Y=135760
X335 1 4 sky130_fd_sc_hd__diode_2 $T=143520 127840 0 0 $X=143330 $Y=127600
X336 1 62 sky130_fd_sc_hd__diode_2 $T=146280 149600 1 0 $X=146090 $Y=146640
X337 1 76 sky130_fd_sc_hd__diode_2 $T=161460 127840 1 0 $X=161270 $Y=124880
X338 1 79 sky130_fd_sc_hd__diode_2 $T=162380 133280 1 0 $X=162190 $Y=130320
X339 1 355 sky130_fd_sc_hd__diode_2 $T=166520 138720 1 0 $X=166330 $Y=135760
X340 1 83 sky130_fd_sc_hd__diode_2 $T=169740 149600 1 0 $X=169550 $Y=146640
X341 1 359 sky130_fd_sc_hd__diode_2 $T=173420 144160 1 0 $X=173230 $Y=141200
X342 1 4 sky130_fd_sc_hd__diode_2 $T=175260 133280 0 0 $X=175070 $Y=133040
X343 1 88 sky130_fd_sc_hd__diode_2 $T=189980 138720 0 0 $X=189790 $Y=138480
X344 1 90 sky130_fd_sc_hd__diode_2 $T=191360 149600 1 0 $X=191170 $Y=146640
X345 1 89 sky130_fd_sc_hd__diode_2 $T=191820 133280 0 0 $X=191630 $Y=133040
X346 1 361 sky130_fd_sc_hd__diode_2 $T=193200 144160 1 0 $X=193010 $Y=141200
X347 1 93 sky130_fd_sc_hd__diode_2 $T=195040 138720 1 0 $X=194850 $Y=135760
X348 1 94 sky130_fd_sc_hd__diode_2 $T=196880 133280 0 0 $X=196690 $Y=133040
X349 1 4 sky130_fd_sc_hd__diode_2 $T=207000 144160 0 0 $X=206810 $Y=143920
X350 1 105 sky130_fd_sc_hd__diode_2 $T=209760 138720 0 0 $X=209570 $Y=138480
X351 1 66 sky130_fd_sc_hd__diode_2 $T=217580 138720 0 0 $X=217390 $Y=138480
X352 1 91 sky130_fd_sc_hd__diode_2 $T=222180 127840 0 0 $X=221990 $Y=127600
X353 1 110 sky130_fd_sc_hd__diode_2 $T=222640 144160 1 0 $X=222450 $Y=141200
X354 1 114 sky130_fd_sc_hd__diode_2 $T=227240 127840 1 0 $X=227050 $Y=124880
X355 1 99 sky130_fd_sc_hd__diode_2 $T=228160 133280 1 0 $X=227970 $Y=130320
X356 1 115 sky130_fd_sc_hd__diode_2 $T=231380 138720 0 0 $X=231190 $Y=138480
X357 1 122 sky130_fd_sc_hd__diode_2 $T=236440 138720 1 0 $X=236250 $Y=135760
X358 1 108 sky130_fd_sc_hd__diode_2 $T=237360 127840 1 0 $X=237170 $Y=124880
X359 1 121 sky130_fd_sc_hd__diode_2 $T=237820 127840 0 0 $X=237630 $Y=127600
X360 1 124 sky130_fd_sc_hd__diode_2 $T=240120 138720 1 0 $X=239930 $Y=135760
X361 1 125 sky130_fd_sc_hd__diode_2 $T=247480 127840 1 0 $X=247290 $Y=124880
X362 1 110 sky130_fd_sc_hd__diode_2 $T=251620 127840 1 0 $X=251430 $Y=124880
X363 1 127 sky130_fd_sc_hd__diode_2 $T=256220 149600 1 0 $X=256030 $Y=146640
X364 1 38 sky130_fd_sc_hd__diode_2 $T=259440 127840 0 0 $X=259250 $Y=127600
X365 1 374 sky130_fd_sc_hd__diode_2 $T=259440 138720 0 0 $X=259250 $Y=138480
X366 1 4 sky130_fd_sc_hd__diode_2 $T=260360 149600 1 0 $X=260170 $Y=146640
X367 1 381 sky130_fd_sc_hd__diode_2 $T=276000 149600 1 0 $X=275810 $Y=146640
X368 1 136 sky130_fd_sc_hd__diode_2 $T=276460 144160 0 0 $X=276270 $Y=143920
X369 1 139 sky130_fd_sc_hd__diode_2 $T=283820 149600 1 0 $X=283630 $Y=146640
X370 1 4 sky130_fd_sc_hd__diode_2 $T=289800 127840 0 0 $X=289610 $Y=127600
X371 1 149 sky130_fd_sc_hd__diode_2 $T=294400 133280 0 0 $X=294210 $Y=133040
X372 1 141 sky130_fd_sc_hd__diode_2 $T=294860 144160 0 0 $X=294670 $Y=143920
X373 1 150 sky130_fd_sc_hd__diode_2 $T=301300 133280 0 0 $X=301110 $Y=133040
X374 1 156 sky130_fd_sc_hd__diode_2 $T=301760 138720 0 0 $X=301570 $Y=138480
X375 1 150 sky130_fd_sc_hd__diode_2 $T=306360 149600 1 0 $X=306170 $Y=146640
X376 1 155 sky130_fd_sc_hd__diode_2 $T=308660 133280 0 0 $X=308470 $Y=133040
X377 1 388 sky130_fd_sc_hd__diode_2 $T=310960 138720 1 0 $X=310770 $Y=135760
X378 1 389 sky130_fd_sc_hd__diode_2 $T=324300 138720 0 0 $X=324110 $Y=138480
X379 1 167 sky130_fd_sc_hd__diode_2 $T=325220 133280 0 0 $X=325030 $Y=133040
X380 1 168 sky130_fd_sc_hd__diode_2 $T=329360 144160 0 0 $X=329170 $Y=143920
X381 1 171 sky130_fd_sc_hd__diode_2 $T=331200 149600 1 0 $X=331010 $Y=146640
X382 1 85 sky130_fd_sc_hd__diode_2 $T=338100 133280 0 0 $X=337910 $Y=133040
X383 1 16 sky130_fd_sc_hd__diode_2 $T=338560 127840 0 0 $X=338370 $Y=127600
X384 1 172 sky130_fd_sc_hd__diode_2 $T=339940 144160 0 0 $X=339750 $Y=143920
X385 1 2 322 ICV_4 $T=35420 138720 1 0 $X=35230 $Y=135760
X386 1 2 17 ICV_4 $T=41400 133280 0 0 $X=41210 $Y=133040
X387 1 2 20 ICV_4 $T=47840 138720 0 0 $X=47650 $Y=138480
X388 1 2 312 ICV_4 $T=50600 138720 1 0 $X=50410 $Y=135760
X389 1 2 327 ICV_4 $T=51520 127840 0 0 $X=51330 $Y=127600
X390 1 2 28 ICV_4 $T=65780 127840 1 0 $X=65590 $Y=124880
X391 1 2 37 ICV_4 $T=86940 144160 0 0 $X=86750 $Y=143920
X392 1 2 51 ICV_4 $T=115000 149600 1 0 $X=114810 $Y=146640
X393 1 2 58 ICV_4 $T=129260 127840 1 0 $X=129070 $Y=124880
X394 1 2 50 ICV_4 $T=129260 133280 1 0 $X=129070 $Y=130320
X395 1 2 54 ICV_4 $T=138460 144160 1 0 $X=138270 $Y=141200
X396 1 2 69 ICV_4 $T=143060 138720 0 0 $X=142870 $Y=138480
X397 1 2 349 ICV_4 $T=145360 138720 1 0 $X=145170 $Y=135760
X398 1 2 77 ICV_4 $T=171120 133280 0 0 $X=170930 $Y=133040
X399 1 2 357 ICV_4 $T=177100 133280 1 0 $X=176910 $Y=130320
X400 1 2 95 ICV_4 $T=196880 138720 0 0 $X=196690 $Y=138480
X401 1 2 362 ICV_4 $T=199180 138720 1 0 $X=198990 $Y=135760
X402 1 2 362 ICV_4 $T=202400 138720 1 0 $X=202210 $Y=135760
X403 1 2 99 ICV_4 $T=202400 144160 1 0 $X=202210 $Y=141200
X404 1 2 364 ICV_4 $T=211600 138720 1 0 $X=211410 $Y=135760
X405 1 2 26 ICV_4 $T=217120 127840 0 0 $X=216930 $Y=127600
X406 1 2 72 ICV_4 $T=218500 127840 1 0 $X=218310 $Y=124880
X407 1 2 113 ICV_4 $T=226780 138720 0 0 $X=226590 $Y=138480
X408 1 2 108 ICV_4 $T=227240 138720 1 0 $X=227050 $Y=135760
X409 1 2 115 ICV_4 $T=237360 133280 0 0 $X=237170 $Y=133040
X410 1 2 4 ICV_4 $T=255300 133280 0 0 $X=255110 $Y=133040
X411 1 2 128 ICV_4 $T=258520 133280 1 0 $X=258330 $Y=130320
X412 1 2 142 ICV_4 $T=286580 127840 1 0 $X=286390 $Y=124880
X413 1 2 151 ICV_4 $T=297620 144160 1 0 $X=297430 $Y=141200
X414 1 2 155 ICV_4 $T=304060 144160 0 0 $X=303870 $Y=143920
X415 1 2 98 ICV_4 $T=305440 138720 1 0 $X=305250 $Y=135760
X416 1 2 159 ICV_4 $T=310960 138720 0 0 $X=310770 $Y=138480
X417 1 2 309 ICV_4 $T=314640 144160 1 0 $X=314450 $Y=141200
X418 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=14720 133280 1 0 $X=14530 $Y=130320
X419 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=27140 138720 0 0 $X=26950 $Y=138480
X420 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=53820 127840 1 0 $X=53630 $Y=124880
X421 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58420 138720 0 0 $X=58230 $Y=138480
X422 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=62100 127840 0 0 $X=61910 $Y=127600
X423 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 127840 0 0 $X=89970 $Y=127600
X424 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 133280 0 0 $X=89970 $Y=133040
X425 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=92460 127840 1 0 $X=92270 $Y=124880
X426 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101200 149600 1 0 $X=101010 $Y=146640
X427 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 127840 1 0 $X=114810 $Y=124880
X428 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=118220 144160 0 0 $X=118030 $Y=143920
X429 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=119140 149600 1 0 $X=118950 $Y=146640
X430 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129260 144160 1 0 $X=129070 $Y=141200
X431 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129260 149600 1 0 $X=129070 $Y=146640
X432 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 133280 1 0 $X=132290 $Y=130320
X433 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=139380 144160 0 0 $X=139190 $Y=143920
X434 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=140300 127840 0 0 $X=140110 $Y=127600
X435 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=147660 127840 1 0 $X=147470 $Y=124880
X436 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=156860 144160 1 0 $X=156670 $Y=141200
X437 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=166980 144160 1 0 $X=166790 $Y=141200
X438 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 149600 1 0 $X=185190 $Y=146640
X439 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=188600 138720 1 0 $X=188410 $Y=135760
X440 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=188600 149600 1 0 $X=188410 $Y=146640
X441 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213440 133280 0 0 $X=213250 $Y=133040
X442 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 133280 1 0 $X=216470 $Y=130320
X443 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=223100 127840 0 0 $X=222910 $Y=127600
X444 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=237360 138720 1 0 $X=237170 $Y=135760
X445 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241040 138720 1 0 $X=240850 $Y=135760
X446 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244260 133280 0 0 $X=244070 $Y=133040
X447 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 127840 1 0 $X=244530 $Y=124880
X448 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 138720 1 0 $X=244530 $Y=135760
X449 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=248400 127840 1 0 $X=248210 $Y=124880
X450 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=250240 144160 1 0 $X=250050 $Y=141200
X451 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=257140 149600 1 0 $X=256950 $Y=146640
X452 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=261280 149600 1 0 $X=261090 $Y=146640
X453 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269100 144160 1 0 $X=268910 $Y=141200
X454 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=271400 127840 0 0 $X=271210 $Y=127600
X455 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=272780 149600 1 0 $X=272590 $Y=146640
X456 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=273240 133280 0 0 $X=273050 $Y=133040
X457 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=279220 138720 0 0 $X=279030 $Y=138480
X458 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=286580 127840 0 0 $X=286390 $Y=127600
X459 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=291640 133280 0 0 $X=291450 $Y=133040
X460 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=303140 149600 1 0 $X=302950 $Y=146640
X461 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 127840 0 0 $X=314450 $Y=127600
X462 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331200 133280 0 0 $X=331010 $Y=133040
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331660 127840 0 0 $X=331470 $Y=127600
X464 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=332120 149600 1 0 $X=331930 $Y=146640
X465 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339020 133280 0 0 $X=338830 $Y=133040
X466 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 127840 0 0 $X=339290 $Y=127600
X467 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=345920 144160 1 0 $X=345730 $Y=141200
X468 1 3 4 ICV_7 $T=7820 138720 1 0 $X=7630 $Y=135760
X469 1 3 311 ICV_7 $T=7820 144160 1 0 $X=7630 $Y=141200
X470 1 316 8 ICV_7 $T=24380 133280 0 0 $X=24190 $Y=133040
X471 1 8 317 ICV_7 $T=25300 127840 1 0 $X=25110 $Y=124880
X472 1 319 312 ICV_7 $T=27600 144160 0 0 $X=27410 $Y=143920
X473 1 9 322 ICV_7 $T=28060 133280 0 0 $X=27870 $Y=133040
X474 1 321 12 ICV_7 $T=29900 127840 0 0 $X=29710 $Y=127600
X475 1 316 14 ICV_7 $T=29900 138720 0 0 $X=29710 $Y=138480
X476 1 15 16 ICV_7 $T=34040 127840 1 0 $X=33850 $Y=124880
X477 1 324 317 ICV_7 $T=34500 133280 1 0 $X=34310 $Y=130320
X478 1 324 322 ICV_7 $T=38180 133280 1 0 $X=37990 $Y=130320
X479 1 326 327 ICV_7 $T=44160 133280 0 0 $X=43970 $Y=133040
X480 1 312 329 ICV_7 $T=44160 144160 1 0 $X=43970 $Y=141200
X481 1 9 22 ICV_7 $T=47840 133280 0 0 $X=47650 $Y=133040
X482 1 8 322 ICV_7 $T=50600 133280 1 0 $X=50410 $Y=130320
X483 1 4 331 ICV_7 $T=54280 127840 0 0 $X=54090 $Y=127600
X484 1 8 330 ICV_7 $T=55660 138720 0 0 $X=55470 $Y=138480
X485 1 4 332 ICV_7 $T=63020 138720 0 0 $X=62830 $Y=138480
X486 1 338 339 ICV_7 $T=79120 138720 0 0 $X=78930 $Y=138480
X487 1 340 55 ICV_7 $T=119140 133280 0 0 $X=118950 $Y=133040
X488 1 33 35 ICV_7 $T=120520 138720 0 0 $X=120330 $Y=138480
X489 1 342 62 ICV_7 $T=126500 144160 1 0 $X=126310 $Y=141200
X490 1 65 67 ICV_7 $T=134320 138720 0 0 $X=134130 $Y=138480
X491 1 344 35 ICV_7 $T=136160 133280 0 0 $X=135970 $Y=133040
X492 1 54 346 ICV_7 $T=137540 127840 0 0 $X=137350 $Y=127600
X493 1 33 347 ICV_7 $T=139840 133280 0 0 $X=139650 $Y=133040
X494 1 67 66 ICV_7 $T=142140 144160 0 0 $X=141950 $Y=143920
X495 1 349 70 ICV_7 $T=148580 144160 1 0 $X=148390 $Y=141200
X496 1 350 70 ICV_7 $T=149500 138720 0 0 $X=149310 $Y=138480
X497 1 62 71 ICV_7 $T=154560 133280 0 0 $X=154370 $Y=133040
X498 1 351 74 ICV_7 $T=158700 138720 0 0 $X=158510 $Y=138480
X499 1 351 75 ICV_7 $T=158700 144160 0 0 $X=158510 $Y=143920
X500 1 80 77 ICV_7 $T=162380 138720 0 0 $X=162190 $Y=138480
X501 1 78 352 ICV_7 $T=162380 149600 1 0 $X=162190 $Y=146640
X502 1 4 354 ICV_7 $T=164220 127840 0 0 $X=164030 $Y=127600
X503 1 358 78 ICV_7 $T=169740 144160 1 0 $X=169550 $Y=141200
X504 1 75 75 ICV_7 $T=170200 144160 0 0 $X=170010 $Y=143920
X505 1 4 96 ICV_7 $T=195960 144160 0 0 $X=195770 $Y=143920
X506 1 101 104 ICV_7 $T=204700 127840 1 0 $X=204510 $Y=124880
X507 1 108 365 ICV_7 $T=216200 133280 0 0 $X=216010 $Y=133040
X508 1 4 367 ICV_7 $T=220340 144160 0 0 $X=220150 $Y=143920
X509 1 91 113 ICV_7 $T=222180 133280 0 0 $X=221990 $Y=133040
X510 1 368 4 ICV_7 $T=226320 127840 0 0 $X=226130 $Y=127600
X511 1 110 61 ICV_7 $T=226320 133280 0 0 $X=226130 $Y=133040
X512 1 105 373 ICV_7 $T=247480 133280 0 0 $X=247290 $Y=133040
X513 1 376 377 ICV_7 $T=251620 133280 0 0 $X=251430 $Y=133040
X514 1 378 379 ICV_7 $T=254380 127840 0 0 $X=254190 $Y=127600
X515 1 109 128 ICV_7 $T=262660 127840 1 0 $X=262470 $Y=124880
X516 1 131 379 ICV_7 $T=268640 127840 0 0 $X=268450 $Y=127600
X517 1 380 136 ICV_7 $T=272780 144160 0 0 $X=272590 $Y=143920
X518 1 131 135 ICV_7 $T=274160 127840 0 0 $X=273970 $Y=127600
X519 1 4 382 ICV_7 $T=276460 133280 0 0 $X=276270 $Y=133040
X520 1 4 383 ICV_7 $T=276460 138720 0 0 $X=276270 $Y=138480
X521 1 137 140 ICV_7 $T=282440 138720 0 0 $X=282250 $Y=138480
X522 1 146 385 ICV_7 $T=292560 138720 0 0 $X=292370 $Y=138480
X523 1 148 144 ICV_7 $T=293020 149600 1 0 $X=292830 $Y=146640
X524 1 139 152 ICV_7 $T=296700 149600 1 0 $X=296510 $Y=146640
X525 1 154 153 ICV_7 $T=301760 144160 1 0 $X=301570 $Y=141200
X526 1 161 387 ICV_7 $T=310040 127840 0 0 $X=309850 $Y=127600
X527 1 161 390 ICV_7 $T=316020 133280 0 0 $X=315830 $Y=133040
X528 1 4 162 ICV_7 $T=316940 127840 1 0 $X=316750 $Y=124880
X529 1 165 4 ICV_7 $T=317400 127840 0 0 $X=317210 $Y=127600
X530 1 158 157 ICV_7 $T=320620 138720 0 0 $X=320430 $Y=138480
X531 1 157 166 ICV_7 $T=321080 149600 1 0 $X=320890 $Y=146640
X532 1 4 169 ICV_7 $T=328900 138720 0 0 $X=328710 $Y=138480
X533 1 3 4 ICV_7 $T=334420 133280 0 0 $X=334230 $Y=133040
X534 1 3 4 ICV_7 $T=334880 127840 0 0 $X=334690 $Y=127600
X535 1 3 4 ICV_7 $T=336260 144160 0 0 $X=336070 $Y=143920
X536 1 2 3 309 4 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 138720 0 0 $X=7630 $Y=138480
X537 1 2 3 311 4 2 6 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 144160 0 0 $X=7630 $Y=143920
X538 1 2 393 310 4 2 7 1 sky130_fd_sc_hd__dfrtp_4 $T=8280 127840 0 0 $X=8090 $Y=127600
X539 1 2 394 314 4 2 311 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 144160 1 0 $X=20970 $Y=141200
X540 1 2 395 323 4 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 144160 0 0 $X=34770 $Y=143920
X541 1 2 396 331 4 2 27 1 sky130_fd_sc_hd__dfrtp_4 $T=54280 133280 1 0 $X=54090 $Y=130320
X542 1 2 397 332 4 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=61640 144160 1 0 $X=61450 $Y=141200
X543 1 2 398 334 4 2 36 1 sky130_fd_sc_hd__dfrtp_4 $T=70380 133280 0 0 $X=70190 $Y=133040
X544 1 2 399 40 4 2 45 1 sky130_fd_sc_hd__dfrtp_4 $T=95220 127840 0 0 $X=95030 $Y=127600
X545 1 2 400 41 4 2 46 1 sky130_fd_sc_hd__dfrtp_4 $T=95220 133280 0 0 $X=95030 $Y=133040
X546 1 2 401 42 4 2 48 1 sky130_fd_sc_hd__dfrtp_4 $T=97980 144160 0 0 $X=97790 $Y=143920
X547 1 2 402 43 4 2 47 1 sky130_fd_sc_hd__dfrtp_4 $T=105340 133280 1 0 $X=105150 $Y=130320
X548 1 2 403 340 4 2 55 1 sky130_fd_sc_hd__dfrtp_4 $T=115920 138720 1 0 $X=115730 $Y=135760
X549 1 2 404 52 4 2 63 1 sky130_fd_sc_hd__dfrtp_4 $T=119140 127840 0 0 $X=118950 $Y=127600
X550 1 2 405 348 4 2 71 1 sky130_fd_sc_hd__dfrtp_4 $T=143520 133280 1 0 $X=143330 $Y=130320
X551 1 2 406 354 4 2 79 1 sky130_fd_sc_hd__dfrtp_4 $T=164220 133280 1 0 $X=164030 $Y=130320
X552 1 2 407 357 4 2 87 1 sky130_fd_sc_hd__dfrtp_4 $T=177100 133280 0 0 $X=176910 $Y=133040
X553 1 2 408 360 4 2 88 1 sky130_fd_sc_hd__dfrtp_4 $T=177560 138720 0 0 $X=177370 $Y=138480
X554 1 2 409 92 4 2 100 1 sky130_fd_sc_hd__dfrtp_4 $T=193200 127840 1 0 $X=193010 $Y=124880
X555 1 2 410 96 4 2 103 1 sky130_fd_sc_hd__dfrtp_4 $T=195960 149600 1 0 $X=195770 $Y=146640
X556 1 2 411 363 4 2 107 1 sky130_fd_sc_hd__dfrtp_4 $T=208840 144160 0 0 $X=208650 $Y=143920
X557 1 2 412 367 4 2 116 1 sky130_fd_sc_hd__dfrtp_4 $T=218960 149600 1 0 $X=218770 $Y=146640
X558 1 2 413 368 4 2 122 1 sky130_fd_sc_hd__dfrtp_4 $T=230000 133280 1 0 $X=229810 $Y=130320
X559 1 2 414 372 4 2 124 1 sky130_fd_sc_hd__dfrtp_4 $T=235520 138720 0 0 $X=235330 $Y=138480
X560 1 2 415 375 4 2 126 1 sky130_fd_sc_hd__dfrtp_4 $T=253000 144160 1 0 $X=252810 $Y=141200
X561 1 2 416 377 4 2 130 1 sky130_fd_sc_hd__dfrtp_4 $T=255300 138720 1 0 $X=255110 $Y=135760
X562 1 2 417 382 4 2 138 1 sky130_fd_sc_hd__dfrtp_4 $T=276460 138720 1 0 $X=276270 $Y=135760
X563 1 2 418 383 4 2 137 1 sky130_fd_sc_hd__dfrtp_4 $T=276460 144160 1 0 $X=276270 $Y=141200
X564 1 2 419 384 4 2 149 1 sky130_fd_sc_hd__dfrtp_4 $T=291640 127840 0 0 $X=291450 $Y=127600
X565 1 2 420 160 4 2 309 1 sky130_fd_sc_hd__dfrtp_4 $T=308200 149600 1 0 $X=308010 $Y=146640
X566 1 2 421 391 4 2 167 1 sky130_fd_sc_hd__dfrtp_4 $T=321080 127840 0 0 $X=320890 $Y=127600
X567 1 2 422 169 4 2 168 1 sky130_fd_sc_hd__dfrtp_4 $T=329820 144160 1 0 $X=329630 $Y=141200
X568 1 2 3 88 4 2 173 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 127840 1 0 $X=334230 $Y=124880
X569 1 2 3 85 4 2 174 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 138720 1 0 $X=334230 $Y=135760
X570 1 2 3 16 4 2 175 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 133280 1 0 $X=334690 $Y=130320
X571 1 2 3 172 4 2 176 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 149600 1 0 $X=334690 $Y=146640
X572 1 313 ICV_15 $T=17940 133280 1 0 $X=17750 $Y=130320
X573 1 13 ICV_15 $T=31740 133280 0 0 $X=31550 $Y=133040
X574 1 328 ICV_15 $T=46000 138720 1 0 $X=45810 $Y=135760
X575 1 26 ICV_15 $T=59800 133280 0 0 $X=59610 $Y=133040
X576 1 335 ICV_15 $T=74060 144160 1 0 $X=73870 $Y=141200
X577 1 38 ICV_15 $T=87860 138720 0 0 $X=87670 $Y=138480
X578 1 4 ICV_15 $T=102120 127840 1 0 $X=101930 $Y=124880
X579 1 43 ICV_15 $T=102120 133280 1 0 $X=101930 $Y=130320
X580 1 4 ICV_15 $T=115920 127840 0 0 $X=115730 $Y=127600
X581 1 4 ICV_15 $T=115920 133280 0 0 $X=115730 $Y=133040
X582 1 359 ICV_15 $T=172040 138720 0 0 $X=171850 $Y=138480
X583 1 20 ICV_15 $T=200100 127840 0 0 $X=199910 $Y=127600
X584 1 98 ICV_15 $T=200100 138720 0 0 $X=199910 $Y=138480
X585 1 106 ICV_15 $T=214360 127840 1 0 $X=214170 $Y=124880
X586 1 107 ICV_15 $T=214360 138720 1 0 $X=214170 $Y=135760
X587 1 126 ICV_15 $T=256220 144160 0 0 $X=256030 $Y=143920
X588 1 141 ICV_15 $T=284280 144160 0 0 $X=284090 $Y=143920
X589 1 2 309 ICV_16 $T=7820 133280 0 0 $X=7630 $Y=133040
X590 1 2 4 ICV_16 $T=7820 149600 1 0 $X=7630 $Y=146640
X591 1 2 4 ICV_16 $T=8280 127840 1 0 $X=8090 $Y=124880
X592 1 2 310 ICV_16 $T=8280 133280 1 0 $X=8090 $Y=130320
X593 1 2 23 ICV_16 $T=55200 144160 0 0 $X=55010 $Y=143920
X594 1 2 27 ICV_16 $T=65320 138720 1 0 $X=65130 $Y=135760
X595 1 2 333 ICV_16 $T=68540 149600 1 0 $X=68350 $Y=146640
X596 1 2 24 ICV_16 $T=71300 127840 0 0 $X=71110 $Y=127600
X597 1 2 36 ICV_16 $T=81880 133280 0 0 $X=81690 $Y=133040
X598 1 2 39 ICV_16 $T=90160 138720 1 0 $X=89970 $Y=135760
X599 1 2 339 ICV_16 $T=90160 144160 1 0 $X=89970 $Y=141200
X600 1 2 40 ICV_16 $T=95220 127840 1 0 $X=95030 $Y=124880
X601 1 2 41 ICV_16 $T=95220 133280 1 0 $X=95030 $Y=130320
X602 1 2 52 ICV_16 $T=118220 127840 1 0 $X=118030 $Y=124880
X603 1 2 348 ICV_16 $T=147200 127840 0 0 $X=147010 $Y=127600
X604 1 2 72 ICV_16 $T=155940 127840 0 0 $X=155750 $Y=127600
X605 1 2 86 ICV_16 $T=178940 149600 1 0 $X=178750 $Y=146640
X606 1 2 87 ICV_16 $T=180320 133280 1 0 $X=180130 $Y=130320
X607 1 2 80 ICV_16 $T=181700 144160 1 0 $X=181510 $Y=141200
X608 1 2 78 ICV_16 $T=182620 144160 0 0 $X=182430 $Y=143920
X609 1 2 100 ICV_16 $T=202400 133280 1 0 $X=202210 $Y=130320
X610 1 2 103 ICV_16 $T=205160 138720 1 0 $X=204970 $Y=135760
X611 1 2 363 ICV_16 $T=208840 149600 1 0 $X=208650 $Y=146640
X612 1 2 366 ICV_16 $T=219880 133280 1 0 $X=219690 $Y=130320
X613 1 2 370 ICV_16 $T=230460 149600 1 0 $X=230270 $Y=146640
X614 1 2 372 ICV_16 $T=235520 144160 1 0 $X=235330 $Y=141200
X615 1 2 133 ICV_16 $T=265420 144160 0 0 $X=265230 $Y=143920
X616 1 2 130 ICV_16 $T=266340 138720 0 0 $X=266150 $Y=138480
X617 1 2 131 ICV_16 $T=266800 133280 0 0 $X=266610 $Y=133040
X618 1 2 143 ICV_16 $T=287960 138720 1 0 $X=287770 $Y=135760
X619 1 2 384 ICV_16 $T=291640 133280 1 0 $X=291450 $Y=130320
X620 1 2 391 ICV_16 $T=321080 127840 1 0 $X=320890 $Y=124880
X621 1 2 392 ICV_16 $T=321080 138720 1 0 $X=320890 $Y=135760
X622 1 2 311 2 316 1 sky130_fd_sc_hd__inv_8 $T=21620 144160 0 0 $X=21430 $Y=143920
X623 1 2 7 2 317 1 sky130_fd_sc_hd__inv_8 $T=22540 127840 0 0 $X=22350 $Y=127600
X624 1 2 18 2 324 1 sky130_fd_sc_hd__inv_8 $T=39100 144160 1 0 $X=38910 $Y=141200
X625 1 2 23 2 328 1 sky130_fd_sc_hd__inv_8 $T=53820 149600 1 0 $X=53630 $Y=146640
X626 1 2 27 2 327 1 sky130_fd_sc_hd__inv_8 $T=63020 133280 0 0 $X=62830 $Y=133040
X627 1 2 32 2 336 1 sky130_fd_sc_hd__inv_8 $T=73140 138720 0 0 $X=72950 $Y=138480
X628 1 2 34 2 29 1 sky130_fd_sc_hd__inv_8 $T=77280 127840 1 0 $X=77090 $Y=124880
X629 1 2 36 2 339 1 sky130_fd_sc_hd__inv_8 $T=80960 138720 1 0 $X=80770 $Y=135760
X630 1 2 45 2 44 1 sky130_fd_sc_hd__inv_8 $T=105340 127840 1 0 $X=105150 $Y=124880
X631 1 2 46 2 49 1 sky130_fd_sc_hd__inv_8 $T=109480 127840 0 0 $X=109290 $Y=127600
X632 1 2 47 2 50 1 sky130_fd_sc_hd__inv_8 $T=109480 133280 0 0 $X=109290 $Y=133040
X633 1 2 57 2 56 1 sky130_fd_sc_hd__inv_8 $T=121900 149600 1 0 $X=121710 $Y=146640
X634 1 2 55 2 342 1 sky130_fd_sc_hd__inv_8 $T=122820 133280 0 0 $X=122630 $Y=133040
X635 1 2 63 2 64 1 sky130_fd_sc_hd__inv_8 $T=132480 127840 0 0 $X=132290 $Y=127600
X636 1 2 71 2 349 1 sky130_fd_sc_hd__inv_8 $T=149500 133280 0 0 $X=149310 $Y=133040
X637 1 2 73 2 347 1 sky130_fd_sc_hd__inv_8 $T=150880 127840 1 0 $X=150690 $Y=124880
X638 1 2 79 2 351 1 sky130_fd_sc_hd__inv_8 $T=166060 133280 0 0 $X=165870 $Y=133040
X639 1 2 85 2 76 1 sky130_fd_sc_hd__inv_8 $T=173880 127840 1 0 $X=173690 $Y=124880
X640 1 2 87 2 83 1 sky130_fd_sc_hd__inv_8 $T=180320 138720 1 0 $X=180130 $Y=135760
X641 1 2 88 2 359 1 sky130_fd_sc_hd__inv_8 $T=191820 138720 0 0 $X=191630 $Y=138480
X642 1 2 100 2 102 1 sky130_fd_sc_hd__inv_8 $T=203320 127840 0 0 $X=203130 $Y=127600
X643 1 2 103 2 362 1 sky130_fd_sc_hd__inv_8 $T=205160 144160 1 0 $X=204970 $Y=141200
X644 1 2 107 2 365 1 sky130_fd_sc_hd__inv_8 $T=217580 144160 1 0 $X=217390 $Y=141200
X645 1 2 122 2 119 1 sky130_fd_sc_hd__inv_8 $T=232300 133280 0 0 $X=232110 $Y=133040
X646 1 2 124 2 114 1 sky130_fd_sc_hd__inv_8 $T=240120 133280 0 0 $X=239930 $Y=133040
X647 1 2 126 2 374 1 sky130_fd_sc_hd__inv_8 $T=260360 144160 0 0 $X=260170 $Y=143920
X648 1 2 130 2 379 1 sky130_fd_sc_hd__inv_8 $T=261280 138720 0 0 $X=261090 $Y=138480
X649 1 2 133 2 132 1 sky130_fd_sc_hd__inv_8 $T=264500 149600 1 0 $X=264310 $Y=146640
X650 1 2 138 2 144 1 sky130_fd_sc_hd__inv_8 $T=287500 133280 0 0 $X=287310 $Y=133040
X651 1 2 137 2 140 1 sky130_fd_sc_hd__inv_8 $T=287500 138720 0 0 $X=287310 $Y=138480
X652 1 2 147 2 134 1 sky130_fd_sc_hd__inv_8 $T=289800 127840 1 0 $X=289610 $Y=124880
X653 1 2 149 2 151 1 sky130_fd_sc_hd__inv_8 $T=296240 133280 0 0 $X=296050 $Y=133040
X654 1 2 309 2 163 1 sky130_fd_sc_hd__inv_8 $T=315560 138720 0 0 $X=315370 $Y=138480
X655 1 2 165 2 386 1 sky130_fd_sc_hd__inv_8 $T=318780 133280 1 0 $X=318590 $Y=130320
X656 1 2 167 2 392 1 sky130_fd_sc_hd__inv_8 $T=327060 133280 0 0 $X=326870 $Y=133040
X657 1 2 168 2 170 1 sky130_fd_sc_hd__inv_8 $T=331200 144160 0 0 $X=331010 $Y=143920
X658 1 2 312 313 2 310 1 sky130_fd_sc_hd__nor2_4 $T=17940 133280 0 0 $X=17750 $Y=133040
X659 1 2 312 315 2 314 1 sky130_fd_sc_hd__nor2_4 $T=21160 138720 0 0 $X=20970 $Y=138480
X660 1 2 312 319 2 323 1 sky130_fd_sc_hd__nor2_4 $T=29440 149600 1 0 $X=29250 $Y=146640
X661 1 2 312 325 2 19 1 sky130_fd_sc_hd__nor2_4 $T=40020 149600 1 0 $X=39830 $Y=146640
X662 1 2 312 330 2 331 1 sky130_fd_sc_hd__nor2_4 $T=50600 138720 0 0 $X=50410 $Y=138480
X663 1 2 30 333 2 332 1 sky130_fd_sc_hd__nor2_4 $T=68540 144160 0 0 $X=68350 $Y=143920
X664 1 2 30 335 2 334 1 sky130_fd_sc_hd__nor2_4 $T=77280 149600 1 0 $X=77090 $Y=146640
X665 1 2 54 341 2 340 1 sky130_fd_sc_hd__nor2_4 $T=121440 144160 1 0 $X=121250 $Y=141200
X666 1 2 54 346 2 68 1 sky130_fd_sc_hd__nor2_4 $T=135700 133280 1 0 $X=135510 $Y=130320
X667 1 2 54 345 2 348 1 sky130_fd_sc_hd__nor2_4 $T=138000 138720 0 0 $X=137810 $Y=138480
X668 1 2 77 353 2 354 1 sky130_fd_sc_hd__nor2_4 $T=161460 138720 1 0 $X=161270 $Y=135760
X669 1 2 77 355 2 357 1 sky130_fd_sc_hd__nor2_4 $T=166060 138720 0 0 $X=165870 $Y=138480
X670 1 2 77 356 2 360 1 sky130_fd_sc_hd__nor2_4 $T=170660 138720 1 0 $X=170470 $Y=135760
X671 1 2 105 364 2 363 1 sky130_fd_sc_hd__nor2_4 $T=211600 138720 0 0 $X=211410 $Y=138480
X672 1 2 111 112 2 368 1 sky130_fd_sc_hd__nor2_4 $T=221260 127840 1 0 $X=221070 $Y=124880
X673 1 2 105 370 2 367 1 sky130_fd_sc_hd__nor2_4 $T=231380 144160 0 0 $X=231190 $Y=143920
X674 1 2 123 371 2 372 1 sky130_fd_sc_hd__nor2_4 $T=239660 127840 0 0 $X=239470 $Y=127600
X675 1 2 105 373 2 375 1 sky130_fd_sc_hd__nor2_4 $T=247480 138720 1 0 $X=247290 $Y=135760
X676 1 2 101 129 2 377 1 sky130_fd_sc_hd__nor2_4 $T=257600 127840 1 0 $X=257410 $Y=124880
X677 1 2 136 381 2 383 1 sky130_fd_sc_hd__nor2_4 $T=277840 149600 1 0 $X=277650 $Y=146640
X678 1 2 136 380 2 382 1 sky130_fd_sc_hd__nor2_4 $T=278300 144160 0 0 $X=278110 $Y=143920
X679 1 2 146 385 2 384 1 sky130_fd_sc_hd__nor2_4 $T=292560 144160 1 0 $X=292370 $Y=141200
X680 1 2 161 387 2 162 1 sky130_fd_sc_hd__nor2_4 $T=310040 133280 1 0 $X=309850 $Y=130320
X681 1 2 161 390 2 391 1 sky130_fd_sc_hd__nor2_4 $T=316020 138720 1 0 $X=315830 $Y=135760
X682 1 2 317 8 9 320 2 313 1 sky130_fd_sc_hd__o22a_4 $T=27140 133280 1 0 $X=26950 $Y=130320
X683 1 2 316 8 9 318 2 315 1 sky130_fd_sc_hd__o22a_4 $T=28060 138720 1 0 $X=27870 $Y=135760
X684 1 2 324 15 12 321 2 319 1 sky130_fd_sc_hd__o22a_4 $T=34960 127840 0 0 $X=34770 $Y=127600
X685 1 2 328 8 9 329 2 325 1 sky130_fd_sc_hd__o22a_4 $T=49220 144160 1 0 $X=49030 $Y=141200
X686 1 2 327 8 9 326 2 330 1 sky130_fd_sc_hd__o22a_4 $T=51520 133280 0 0 $X=51330 $Y=133040
X687 1 2 336 33 35 337 2 333 1 sky130_fd_sc_hd__o22a_4 $T=79580 144160 0 0 $X=79390 $Y=143920
X688 1 2 339 33 35 338 2 335 1 sky130_fd_sc_hd__o22a_4 $T=82800 144160 1 0 $X=82610 $Y=141200
X689 1 2 342 33 35 343 2 341 1 sky130_fd_sc_hd__o22a_4 $T=124200 138720 0 0 $X=124010 $Y=138480
X690 1 2 347 33 35 344 2 346 1 sky130_fd_sc_hd__o22a_4 $T=138000 138720 1 0 $X=137810 $Y=135760
X691 1 2 349 65 69 350 2 345 1 sky130_fd_sc_hd__o22a_4 $T=141220 144160 1 0 $X=141030 $Y=141200
X692 1 2 351 78 75 352 2 353 1 sky130_fd_sc_hd__o22a_4 $T=162380 144160 0 0 $X=162190 $Y=143920
X693 1 2 359 78 75 358 2 356 1 sky130_fd_sc_hd__o22a_4 $T=171580 149600 1 0 $X=171390 $Y=146640
X694 1 2 83 78 75 86 2 355 1 sky130_fd_sc_hd__o22a_4 $T=175260 144160 0 0 $X=175070 $Y=143920
X695 1 2 362 93 95 361 2 90 1 sky130_fd_sc_hd__o22a_4 $T=195040 144160 1 0 $X=194850 $Y=141200
X696 1 2 365 108 113 366 2 364 1 sky130_fd_sc_hd__o22a_4 $T=219880 138720 1 0 $X=219690 $Y=135760
X697 1 2 115 108 113 369 2 370 1 sky130_fd_sc_hd__o22a_4 $T=226780 144160 1 0 $X=226590 $Y=141200
X698 1 2 114 118 120 117 2 371 1 sky130_fd_sc_hd__o22a_4 $T=229080 127840 1 0 $X=228890 $Y=124880
X699 1 2 374 131 128 376 2 373 1 sky130_fd_sc_hd__o22a_4 $T=259440 133280 0 0 $X=259250 $Y=133040
X700 1 2 379 131 128 378 2 129 1 sky130_fd_sc_hd__o22a_4 $T=261280 127840 0 0 $X=261090 $Y=127600
X701 1 2 140 139 141 145 2 381 1 sky130_fd_sc_hd__o22a_4 $T=285660 149600 1 0 $X=285470 $Y=146640
X702 1 2 144 139 141 143 2 380 1 sky130_fd_sc_hd__o22a_4 $T=287500 144160 0 0 $X=287310 $Y=143920
X703 1 2 151 139 141 154 2 385 1 sky130_fd_sc_hd__o22a_4 $T=296700 144160 0 0 $X=296510 $Y=143920
X704 1 2 386 153 156 388 2 387 1 sky130_fd_sc_hd__o22a_4 $T=303600 138720 0 0 $X=303410 $Y=138480
X705 1 2 392 157 158 389 2 390 1 sky130_fd_sc_hd__o22a_4 $T=317860 144160 1 0 $X=317670 $Y=141200
X706 1 2 10 2 11 1 sky130_fd_sc_hd__buf_1 $T=30820 127840 1 0 $X=30630 $Y=124880
X707 1 2 20 2 322 1 sky130_fd_sc_hd__buf_1 $T=45540 138720 0 0 $X=45350 $Y=138480
X708 1 2 26 2 312 1 sky130_fd_sc_hd__buf_1 $T=63020 138720 1 0 $X=62830 $Y=135760
X709 1 2 67 2 33 1 sky130_fd_sc_hd__buf_1 $T=136160 144160 1 0 $X=135970 $Y=141200
X710 1 2 67 2 65 1 sky130_fd_sc_hd__buf_1 $T=143060 149600 1 0 $X=142870 $Y=146640
X711 1 2 70 2 35 1 sky130_fd_sc_hd__buf_1 $T=147200 138720 0 0 $X=147010 $Y=138480
X712 1 2 70 2 69 1 sky130_fd_sc_hd__buf_1 $T=148120 149600 1 0 $X=147930 $Y=146640
X713 1 2 72 2 8 1 sky130_fd_sc_hd__buf_1 $T=153640 127840 0 0 $X=153450 $Y=127600
X714 1 2 81 2 82 1 sky130_fd_sc_hd__buf_1 $T=166060 127840 1 0 $X=165870 $Y=124880
X715 1 2 89 2 91 1 sky130_fd_sc_hd__buf_1 $T=191820 138720 1 0 $X=191630 $Y=135760
X716 1 2 94 2 20 1 sky130_fd_sc_hd__buf_1 $T=196880 138720 1 0 $X=196690 $Y=135760
X717 1 2 20 2 99 1 sky130_fd_sc_hd__buf_1 $T=200100 133280 1 0 $X=199910 $Y=130320
X718 1 2 97 2 26 1 sky130_fd_sc_hd__buf_1 $T=203320 144160 0 0 $X=203130 $Y=143920
X719 1 2 26 2 101 1 sky130_fd_sc_hd__buf_1 $T=208380 127840 1 0 $X=208190 $Y=124880
X720 1 2 26 2 105 1 sky130_fd_sc_hd__buf_1 $T=214820 127840 0 0 $X=214630 $Y=127600
X721 1 2 91 2 109 1 sky130_fd_sc_hd__buf_1 $T=219880 127840 0 0 $X=219690 $Y=127600
X722 1 2 91 2 110 1 sky130_fd_sc_hd__buf_1 $T=219880 133280 0 0 $X=219690 $Y=133040
X723 1 2 150 2 153 1 sky130_fd_sc_hd__buf_1 $T=298540 138720 0 0 $X=298350 $Y=138480
X724 1 2 150 2 139 1 sky130_fd_sc_hd__buf_1 $T=301760 138720 1 0 $X=301570 $Y=135760
X725 1 2 155 2 156 1 sky130_fd_sc_hd__buf_1 $T=301760 149600 1 0 $X=301570 $Y=146640
X726 1 2 150 2 157 1 sky130_fd_sc_hd__buf_1 $T=307280 144160 0 0 $X=307090 $Y=143920
X727 1 2 155 2 158 1 sky130_fd_sc_hd__buf_1 $T=308660 138720 1 0 $X=308470 $Y=135760
X728 1 2 13 317 322 2 320 1 sky130_fd_sc_hd__o21a_4 $T=34960 133280 0 0 $X=34770 $Y=133040
X729 1 2 14 316 322 2 318 1 sky130_fd_sc_hd__o21a_4 $T=34960 138720 0 0 $X=34770 $Y=138480
X730 1 2 17 324 322 2 321 1 sky130_fd_sc_hd__o21a_4 $T=38180 138720 1 0 $X=37990 $Y=135760
X731 1 2 21 328 322 2 329 1 sky130_fd_sc_hd__o21a_4 $T=48760 144160 0 0 $X=48570 $Y=143920
X732 1 2 22 327 322 2 326 1 sky130_fd_sc_hd__o21a_4 $T=53820 138720 1 0 $X=53630 $Y=135760
X733 1 2 37 336 39 2 337 1 sky130_fd_sc_hd__o21a_4 $T=84640 149600 1 0 $X=84450 $Y=146640
X734 1 2 38 339 39 2 338 1 sky130_fd_sc_hd__o21a_4 $T=91080 138720 0 0 $X=90890 $Y=138480
X735 1 2 59 342 62 2 343 1 sky130_fd_sc_hd__o21a_4 $T=128340 144160 0 0 $X=128150 $Y=143920
X736 1 2 66 349 62 2 350 1 sky130_fd_sc_hd__o21a_4 $T=147200 144160 0 0 $X=147010 $Y=143920
X737 1 2 60 347 62 2 344 1 sky130_fd_sc_hd__o21a_4 $T=148120 138720 1 0 $X=147930 $Y=135760
X738 1 2 74 351 80 2 352 1 sky130_fd_sc_hd__o21a_4 $T=161460 144160 1 0 $X=161270 $Y=141200
X739 1 2 84 359 80 2 358 1 sky130_fd_sc_hd__o21a_4 $T=175260 144160 1 0 $X=175070 $Y=141200
X740 1 2 98 362 99 2 361 1 sky130_fd_sc_hd__o21a_4 $T=203320 138720 0 0 $X=203130 $Y=138480
X741 1 2 66 365 110 2 366 1 sky130_fd_sc_hd__o21a_4 $T=219420 138720 0 0 $X=219230 $Y=138480
X742 1 2 61 115 110 2 369 1 sky130_fd_sc_hd__o21a_4 $T=230000 138720 1 0 $X=229810 $Y=135760
X743 1 2 121 114 99 2 117 1 sky130_fd_sc_hd__o21a_4 $T=231380 127840 0 0 $X=231190 $Y=127600
X744 1 2 59 374 110 2 376 1 sky130_fd_sc_hd__o21a_4 $T=251620 133280 1 0 $X=251430 $Y=130320
X745 1 2 38 379 109 2 378 1 sky130_fd_sc_hd__o21a_4 $T=261740 133280 1 0 $X=261550 $Y=130320
X746 1 2 60 134 109 2 135 1 sky130_fd_sc_hd__o21a_4 $T=273700 127840 1 0 $X=273510 $Y=124880
X747 1 2 98 386 159 2 388 1 sky130_fd_sc_hd__o21a_4 $T=305440 144160 1 0 $X=305250 $Y=141200
X748 1 2 164 392 159 2 389 1 sky130_fd_sc_hd__o21a_4 $T=317860 144160 0 0 $X=317670 $Y=143920
X749 1 2 311 ICV_22 $T=18400 144160 0 0 $X=18210 $Y=143920
X750 1 2 4 ICV_22 $T=30360 144160 0 0 $X=30170 $Y=143920
X751 1 2 9 ICV_22 $T=42320 138720 0 0 $X=42130 $Y=138480
X752 1 2 21 ICV_22 $T=45540 144160 0 0 $X=45350 $Y=143920
X753 1 2 4 ICV_22 $T=67160 133280 0 0 $X=66970 $Y=133040
X754 1 2 42 ICV_22 $T=96600 144160 1 0 $X=96410 $Y=141200
X755 1 2 347 ICV_22 $T=142600 133280 0 0 $X=142410 $Y=133040
X756 1 2 60 ICV_22 $T=146280 133280 0 0 $X=146090 $Y=133040
X757 1 2 356 ICV_22 $T=167440 138720 1 0 $X=167250 $Y=135760
X758 1 2 4 ICV_22 $T=174340 138720 0 0 $X=174150 $Y=138480
X759 1 2 97 ICV_22 $T=198720 144160 0 0 $X=198530 $Y=143920
X760 1 2 365 ICV_22 $T=216660 138720 1 0 $X=216470 $Y=135760
X761 1 2 369 ICV_22 $T=223560 144160 1 0 $X=223370 $Y=141200
X762 1 2 105 ICV_22 $T=226780 144160 0 0 $X=226590 $Y=143920
X763 1 2 4 ICV_22 $T=232300 138720 0 0 $X=232110 $Y=138480
X764 1 2 134 ICV_22 $T=269100 127840 1 0 $X=268910 $Y=124880
X765 1 2 138 ICV_22 $T=282900 133280 0 0 $X=282710 $Y=133040
X766 1 2 150 ICV_22 $T=295320 138720 0 0 $X=295130 $Y=138480
X767 1 2 164 ICV_22 $T=314640 144160 0 0 $X=314450 $Y=143920
X768 1 2 ICV_23 $T=36800 127840 1 0 $X=36610 $Y=124880
X769 1 2 ICV_23 $T=76360 133280 1 0 $X=76170 $Y=130320
X770 1 2 ICV_23 $T=77740 127840 0 0 $X=77550 $Y=127600
X771 1 2 ICV_23 $T=81420 127840 1 0 $X=81230 $Y=124880
X772 1 2 ICV_23 $T=90160 149600 1 0 $X=89970 $Y=146640
X773 1 2 ICV_23 $T=96600 138720 0 0 $X=96410 $Y=138480
X774 1 2 ICV_23 $T=104420 138720 1 0 $X=104230 $Y=135760
X775 1 2 ICV_23 $T=104420 144160 1 0 $X=104230 $Y=141200
X776 1 2 ICV_23 $T=136620 127840 1 0 $X=136430 $Y=124880
X777 1 2 ICV_23 $T=174340 127840 0 0 $X=174150 $Y=127600
X778 1 2 ICV_23 $T=185380 127840 0 0 $X=185190 $Y=127600
X779 1 2 ICV_23 $T=188600 133280 1 0 $X=188410 $Y=130320
X780 1 2 ICV_23 $T=202400 133280 0 0 $X=202210 $Y=133040
X781 1 2 ICV_23 $T=235520 144160 0 0 $X=235330 $Y=143920
X782 1 2 ICV_23 $T=244720 149600 1 0 $X=244530 $Y=146640
X783 1 2 ICV_23 $T=272780 133280 1 0 $X=272590 $Y=130320
X784 1 2 ICV_23 $T=300840 127840 1 0 $X=300650 $Y=124880
X785 1 2 314 312 ICV_27 $T=21160 138720 1 0 $X=20970 $Y=135760
X786 1 2 322 328 ICV_27 $T=49220 149600 1 0 $X=49030 $Y=146640
X787 1 2 33 30 ICV_27 $T=74520 144160 0 0 $X=74330 $Y=143920
X788 1 2 337 35 ICV_27 $T=77740 144160 1 0 $X=77550 $Y=141200
X789 1 2 35 33 ICV_27 $T=82800 138720 0 0 $X=82610 $Y=138480
X790 1 2 39 336 ICV_27 $T=91080 144160 0 0 $X=90890 $Y=143920
X791 1 2 341 57 ICV_27 $T=121440 144160 0 0 $X=121250 $Y=143920
X792 1 2 77 353 ICV_27 $T=161460 133280 0 0 $X=161270 $Y=133040
X793 1 2 84 360 ICV_27 $T=175720 138720 1 0 $X=175530 $Y=135760
X794 1 2 123 371 ICV_27 $T=239660 127840 1 0 $X=239470 $Y=124880
X795 1 2 374 59 ICV_27 $T=249780 127840 0 0 $X=249590 $Y=127600
X796 1 2 4 375 ICV_27 $T=253000 138720 0 0 $X=252810 $Y=138480
X797 1 2 141 139 ICV_27 $T=287960 144160 1 0 $X=287770 $Y=141200
X798 1 2 386 386 ICV_27 $T=303600 133280 0 0 $X=303410 $Y=133040
X799 1 2 4 160 ICV_27 $T=309580 144160 0 0 $X=309390 $Y=143920
X800 1 2 159 392 ICV_27 $T=324300 144160 0 0 $X=324110 $Y=143920
X801 1 2 ICV_29 $T=10580 138720 1 0 $X=10390 $Y=135760
X802 1 2 ICV_29 $T=10580 144160 1 0 $X=10390 $Y=141200
X803 1 2 ICV_29 $T=20240 149600 1 0 $X=20050 $Y=146640
X804 1 2 ICV_29 $T=41400 127840 0 0 $X=41210 $Y=127600
X805 1 2 ICV_29 $T=57960 149600 1 0 $X=57770 $Y=146640
X806 1 2 ICV_29 $T=104420 149600 1 0 $X=104230 $Y=146640
X807 1 2 ICV_29 $T=107640 138720 0 0 $X=107450 $Y=138480
X808 1 2 ICV_29 $T=108560 144160 0 0 $X=108370 $Y=143920
X809 1 2 ICV_29 $T=115920 133280 1 0 $X=115730 $Y=130320
X810 1 2 ICV_29 $T=126960 133280 0 0 $X=126770 $Y=133040
X811 1 2 ICV_29 $T=132480 149600 1 0 $X=132290 $Y=146640
X812 1 2 ICV_29 $T=149500 149600 1 0 $X=149310 $Y=146640
X813 1 2 ICV_29 $T=178020 127840 1 0 $X=177830 $Y=124880
X814 1 2 ICV_29 $T=246560 144160 0 0 $X=246370 $Y=143920
X815 1 2 ICV_29 $T=276920 127840 0 0 $X=276730 $Y=127600
X816 1 2 ICV_29 $T=300840 133280 1 0 $X=300650 $Y=130320
X817 1 2 ICV_29 $T=331660 138720 0 0 $X=331470 $Y=138480
X818 1 2 24 25 2 17 1 sky130_fd_sc_hd__or2_4 $T=57040 127840 1 0 $X=56850 $Y=124880
X819 1 2 24 29 2 13 1 sky130_fd_sc_hd__or2_4 $T=67160 127840 0 0 $X=66970 $Y=127600
X820 1 2 24 31 2 14 1 sky130_fd_sc_hd__or2_4 $T=69000 127840 1 0 $X=68810 $Y=124880
X821 1 2 58 49 2 60 1 sky130_fd_sc_hd__or2_4 $T=125120 127840 1 0 $X=124930 $Y=124880
X822 1 2 58 50 2 61 1 sky130_fd_sc_hd__or2_4 $T=125120 133280 1 0 $X=124930 $Y=130320
X823 1 2 58 64 2 66 1 sky130_fd_sc_hd__or2_4 $T=133400 127840 1 0 $X=133210 $Y=124880
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and2_4 VNB VPB A B VPWR X VGND
** N=38 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 9 A 8 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=760 $Y=235 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1335 $Y=235 $D=9
M3 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1765 $Y=235 $D=9
M4 X 8 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2195 $Y=235 $D=9
M5 VGND 8 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2625 $Y=235 $D=9
M6 8 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M7 VPWR B 8 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1335 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1765 $Y=1485 $D=89
M10 X 8 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2195 $Y=1485 $D=89
M11 VPWR 8 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2625 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor3_4 VNB VPB A B C VPWR Y VGND
** N=63 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=415 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=835 $Y=235 $D=9
M2 Y A VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1255 $Y=235 $D=9
M3 VGND A Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1675 $Y=235 $D=9
M4 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2095 $Y=235 $D=9
M5 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2515 $Y=235 $D=9
M6 Y B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2935 $Y=235 $D=9
M7 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3355 $Y=235 $D=9
M8 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3775 $Y=235 $D=9
M9 VGND C Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4195 $Y=235 $D=9
M10 Y C VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4615 $Y=235 $D=9
M11 VGND B Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5035 $Y=235 $D=9
M12 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=415 $Y=1485 $D=89
M13 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=835 $Y=1485 $D=89
M14 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1255 $Y=1485 $D=89
M15 9 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1675 $Y=1485 $D=89
M16 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2095 $Y=1485 $D=89
M17 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2515 $Y=1485 $D=89
M18 10 B 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2935 $Y=1485 $D=89
M19 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3355 $Y=1485 $D=89
M20 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3775 $Y=1485 $D=89
M21 Y C 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4195 $Y=1485 $D=89
M22 10 C Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4615 $Y=1485 $D=89
M23 9 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5035 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21oi_4 VNB VPB B1 A2 A1 Y VPWR VGND
** N=57 EP=8 IP=0 FDC=24
*.SEEDPROM
M0 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=400 $Y=235 $D=9
M1 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=830 $Y=235 $D=9
M2 Y B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1260 $Y=235 $D=9
M3 VGND B1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1690 $Y=235 $D=9
M4 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2160 $Y=235 $D=9
M5 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2590 $Y=235 $D=9
M6 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3020 $Y=235 $D=9
M7 Y A1 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3450 $Y=235 $D=9
M8 10 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3880 $Y=235 $D=9
M9 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4310 $Y=235 $D=9
M10 10 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4740 $Y=235 $D=9
M11 VGND A2 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5170 $Y=235 $D=9
M12 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M13 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M14 Y B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M15 9 B1 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M16 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2150 $Y=1485 $D=89
M17 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2590 $Y=1485 $D=89
M18 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3020 $Y=1485 $D=89
M19 9 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3450 $Y=1485 $D=89
M20 VPWR A1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3880 $Y=1485 $D=89
M21 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4310 $Y=1485 $D=89
M22 VPWR A2 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4740 $Y=1485 $D=89
M23 9 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_36 1 3 4
** N=4 EP=3 IP=6 FDC=2
*.SEEDPROM
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5 6
** N=6 EP=6 IP=10 FDC=6
*.SEEDPROM
X0 1 3 4 ICV_7 $T=2300 0 0 0 $X=2110 $Y=-240
X1 1 2 5 2 6 1 sky130_fd_sc_hd__buf_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or4_4 VNB VPB D C B A VPWR X VGND
** N=46 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 10 D VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND C 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=950 $Y=235 $D=9
M2 10 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1370 $Y=235 $D=9
M3 VGND A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1790 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2320 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2740 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3160 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3580 $Y=235 $D=9
M8 11 D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M9 12 C 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=950 $Y=1485 $D=88
M10 13 B 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1370 $Y=1485 $D=88
M11 VPWR A 13 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1790 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2320 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2740 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3160 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3580 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and3_4 VNB VPB A B C VPWR X VGND
** N=43 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 10 A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=775 $Y=235 $D=9
M1 11 B 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1320 $Y=235 $D=8
M2 VGND C 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1680 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2255 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2685 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3115 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3545 $Y=235 $D=9
M7 VPWR A 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=775 $Y=1485 $D=89
M8 9 B VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1320 $Y=1485 $D=89
M9 VPWR C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1750 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2255 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2685 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3115 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3545 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__or3_4 VNB VPB C B A VPWR X VGND
** N=49 EP=8 IP=0 FDC=14
*.SEEDPROM
M0 VGND C 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 9 B VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 VGND A 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2185 $Y=235 $D=9
M4 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2605 $Y=235 $D=9
M5 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3025 $Y=235 $D=9
M6 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3445 $Y=235 $D=9
M7 10 C 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M8 11 B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=88
M9 VPWR A 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2185 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2605 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3025 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3445 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4_4 VNB VPB A B C D VPWR X VGND
** N=44 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 11 A 10 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 12 B 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=790 $Y=235 $D=8
M2 13 C 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1275 $Y=235 $D=8
M3 VGND D 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1860 $Y=235 $D=9
M4 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2335 $Y=235 $D=9
M5 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2755 $Y=235 $D=9
M6 X 10 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3175 $Y=235 $D=9
M7 VGND 10 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3595 $Y=235 $D=9
M8 10 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M9 VPWR B 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M10 10 C VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1275 $Y=1485 $D=89
M11 VPWR D 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1855 $Y=1485 $D=89
M12 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2335 $Y=1485 $D=89
M13 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2755 $Y=1485 $D=89
M14 X 10 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3175 $Y=1485 $D=89
M15 VPWR 10 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3595 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21boi_4 VNB VPB B1_N A2 A1 VPWR Y VGND
** N=63 EP=8 IP=0 FDC=26
*.SEEDPROM
M0 VGND B1_N 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=550 $Y=235 $D=9
M1 Y 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1080 $Y=235 $D=9
M2 VGND 9 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1510 $Y=235 $D=9
M3 Y 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1940 $Y=235 $D=9
M4 VGND 9 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2370 $Y=235 $D=9
M5 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3140 $Y=235 $D=9
M6 Y A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3570 $Y=235 $D=9
M7 11 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4000 $Y=235 $D=9
M8 Y A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4430 $Y=235 $D=9
M9 11 A1 Y VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4860 $Y=235 $D=9
M10 VGND A2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5290 $Y=235 $D=9
M11 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5720 $Y=235 $D=9
M12 VGND A2 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6150 $Y=235 $D=9
M13 VPWR B1_N 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=430 $Y=1485 $D=89
M14 Y 9 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1380 $Y=1485 $D=89
M15 10 9 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1810 $Y=1485 $D=89
M16 Y 9 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2240 $Y=1485 $D=89
M17 10 9 Y VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2670 $Y=1485 $D=89
M18 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3130 $Y=1485 $D=89
M19 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3570 $Y=1485 $D=89
M20 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4000 $Y=1485 $D=89
M21 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4430 $Y=1485 $D=89
M22 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4860 $Y=1485 $D=89
M23 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5290 $Y=1485 $D=89
M24 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5720 $Y=1485 $D=89
M25 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6150 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289
** N=788 EP=289 IP=6272 FDC=8453
*.SEEDPROM
M0 1 385 387 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=182295 $Y=95435 $D=9
M1 10 386 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=182725 $Y=95435 $D=9
M2 1 386 10 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=183155 $Y=95435 $D=9
M3 10 386 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=183585 $Y=95435 $D=9
M4 1 386 10 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=184015 $Y=95435 $D=9
M5 386 387 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=184975 $Y=95435 $D=9
M6 1 387 386 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=185395 $Y=95435 $D=9
M7 402 388 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=185855 $Y=95435 $D=9
M8 386 3 402 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=186235 $Y=95435 $D=9
M9 403 3 386 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=186655 $Y=95435 $D=9
M10 1 388 403 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=187075 $Y=95435 $D=9
M11 404 4 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=191755 $Y=83435 $D=9
M12 391 389 404 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=192175 $Y=83435 $D=9
M13 404 389 391 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=192595 $Y=83435 $D=9
M14 1 4 404 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=193015 $Y=83435 $D=9
M15 391 390 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=193435 $Y=83435 $D=9
M16 1 390 391 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=193855 $Y=83435 $D=9
M17 390 5 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=194795 $Y=83435 $D=9
M18 1 6 390 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=195215 $Y=83435 $D=9
M19 390 6 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=195635 $Y=83435 $D=9
M20 1 5 390 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=196055 $Y=83435 $D=9
M21 397 391 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=196475 $Y=83435 $D=9
M22 1 391 397 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=196895 $Y=83435 $D=9
M23 397 391 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=197315 $Y=83435 $D=9
M24 1 391 397 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=197735 $Y=83435 $D=9
M25 1 7 405 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=203715 $Y=100875 $D=9
M26 405 7 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204135 $Y=100875 $D=9
M27 1 8 405 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204555 $Y=100875 $D=9
M28 405 8 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204975 $Y=100875 $D=9
M29 1 9 405 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=205415 $Y=100875 $D=9
M30 405 9 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=205835 $Y=100875 $D=9
M31 405 392 393 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=207275 $Y=100875 $D=9
M32 393 392 405 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=207695 $Y=100875 $D=9
M33 405 3 393 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=208115 $Y=100875 $D=9
M34 393 3 405 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=208565 $Y=100875 $D=9
M35 401 393 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=209505 $Y=100875 $D=9
M36 1 393 401 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=209925 $Y=100875 $D=9
M37 401 393 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=210345 $Y=100875 $D=9
M38 1 393 401 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=210765 $Y=100875 $D=9
M39 2 385 387 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=182295 $Y=96685 $D=89
M40 10 386 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=182725 $Y=96685 $D=89
M41 2 386 10 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=183155 $Y=96685 $D=89
M42 10 386 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=183585 $Y=96685 $D=89
M43 2 386 10 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=184015 $Y=96685 $D=89
M44 386 387 394 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=184975 $Y=96685 $D=89
M45 394 387 386 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=185395 $Y=96685 $D=89
M46 2 388 394 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=185815 $Y=96685 $D=89
M47 394 3 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=186235 $Y=96685 $D=89
M48 2 3 394 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=186655 $Y=96685 $D=89
M49 394 388 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=187075 $Y=96685 $D=89
M50 2 4 395 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=191755 $Y=81835 $D=89
M51 395 389 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=192175 $Y=81835 $D=89
M52 2 389 395 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=192595 $Y=81835 $D=89
M53 395 4 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=193015 $Y=81835 $D=89
M54 391 390 395 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=193435 $Y=81835 $D=89
M55 395 390 391 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=193855 $Y=81835 $D=89
M56 396 5 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=194795 $Y=81835 $D=89
M57 390 6 396 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=195215 $Y=81835 $D=89
M58 396 6 390 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=195635 $Y=81835 $D=89
M59 2 5 396 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=196055 $Y=81835 $D=89
M60 397 391 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=196475 $Y=81835 $D=89
M61 2 391 397 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=196895 $Y=81835 $D=89
M62 397 391 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=197315 $Y=81835 $D=89
M63 2 391 397 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=197735 $Y=81835 $D=89
M64 2 7 398 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=203715 $Y=102125 $D=89
M65 398 7 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204135 $Y=102125 $D=89
M66 399 8 398 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204555 $Y=102125 $D=89
M67 398 8 399 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204975 $Y=102125 $D=89
M68 393 9 399 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=205915 $Y=102125 $D=89
M69 399 9 393 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=206335 $Y=102125 $D=89
M70 2 392 400 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=207275 $Y=102125 $D=89
M71 400 392 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=207695 $Y=102125 $D=89
M72 393 3 400 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=208115 $Y=102125 $D=89
M73 400 3 393 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=208565 $Y=102125 $D=89
M74 401 393 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=209505 $Y=102125 $D=89
M75 2 393 401 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=209925 $Y=102125 $D=89
M76 401 393 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=210345 $Y=102125 $D=89
M77 2 393 401 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=210765 $Y=102125 $D=89
X78 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=80185 $D=191
X79 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=85625 $D=191
X80 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=91065 $D=191
X81 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=96505 $D=191
X82 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=101945 $D=191
X83 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=107385 $D=191
X84 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=112825 $D=191
X85 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=118265 $D=191
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 78880 0 0 $X=5330 $Y=78640
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=10580 95200 1 0 $X=10390 $Y=92240
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28520 106080 1 0 $X=28330 $Y=103120
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=64400 122400 1 0 $X=64210 $Y=119440
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=66700 106080 1 0 $X=66510 $Y=103120
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 84320 0 0 $X=76170 $Y=84080
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=80500 106080 1 0 $X=80310 $Y=103120
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=117300 106080 1 0 $X=117110 $Y=103120
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=137080 95200 1 0 $X=136890 $Y=92240
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=143060 116960 1 0 $X=142870 $Y=114000
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 116960 0 0 $X=144250 $Y=116720
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164220 122400 1 0 $X=164030 $Y=119440
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164680 95200 0 0 $X=164490 $Y=94960
X99 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164680 106080 0 0 $X=164490 $Y=105840
X100 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=188600 100640 1 0 $X=188410 $Y=97680
X101 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 111520 1 0 $X=214630 $Y=108560
X102 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=216660 122400 1 0 $X=216470 $Y=119440
X103 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 116960 0 0 $X=230270 $Y=116720
X104 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=279220 95200 0 0 $X=279030 $Y=94960
X105 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 100640 0 0 $X=284550 $Y=100400
X106 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=288880 84320 1 0 $X=288690 $Y=81360
X107 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=289800 89760 1 0 $X=289610 $Y=86800
X108 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=301760 111520 0 0 $X=301570 $Y=111280
X109 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=304980 106080 1 0 $X=304790 $Y=103120
X110 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=310960 122400 1 0 $X=310770 $Y=119440
X111 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=318320 106080 0 0 $X=318130 $Y=105840
X112 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=347760 106080 1 0 $X=347570 $Y=103120
X113 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 78880 1 180 $X=348950 $Y=78640
X114 1 2 ICV_1 $T=5520 84320 1 0 $X=5330 $Y=81360
X115 1 2 ICV_1 $T=5520 89760 1 0 $X=5330 $Y=86800
X116 1 2 ICV_1 $T=5520 95200 1 0 $X=5330 $Y=92240
X117 1 2 ICV_1 $T=5520 100640 1 0 $X=5330 $Y=97680
X118 1 2 ICV_1 $T=5520 106080 1 0 $X=5330 $Y=103120
X119 1 2 ICV_1 $T=5520 111520 1 0 $X=5330 $Y=108560
X120 1 2 ICV_1 $T=5520 116960 1 0 $X=5330 $Y=114000
X121 1 2 ICV_1 $T=5520 122400 1 0 $X=5330 $Y=119440
X122 1 2 ICV_1 $T=350520 84320 0 180 $X=348950 $Y=81360
X123 1 2 ICV_1 $T=350520 89760 0 180 $X=348950 $Y=86800
X124 1 2 ICV_1 $T=350520 95200 0 180 $X=348950 $Y=92240
X125 1 2 ICV_1 $T=350520 100640 0 180 $X=348950 $Y=97680
X126 1 2 ICV_1 $T=350520 106080 0 180 $X=348950 $Y=103120
X127 1 2 ICV_1 $T=350520 111520 0 180 $X=348950 $Y=108560
X128 1 2 ICV_1 $T=350520 116960 0 180 $X=348950 $Y=114000
X129 1 2 ICV_1 $T=350520 122400 0 180 $X=348950 $Y=119440
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 95200 1 0 $X=6710 $Y=92240
X227 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=10580 100640 1 0 $X=10390 $Y=97680
X228 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=15640 89760 1 0 $X=15450 $Y=86800
X229 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 95200 1 0 $X=15910 $Y=92240
X230 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 106080 1 0 $X=20050 $Y=103120
X231 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 122400 1 0 $X=20050 $Y=119440
X232 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34500 89760 1 0 $X=34310 $Y=86800
X233 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39100 122400 0 0 $X=38910 $Y=122160
X234 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39560 78880 0 0 $X=39370 $Y=78640
X235 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39560 100640 1 0 $X=39370 $Y=97680
X236 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=42780 89760 1 0 $X=42590 $Y=86800
X237 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=43700 122400 1 0 $X=43510 $Y=119440
X238 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=48300 122400 1 0 $X=48110 $Y=119440
X239 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=56580 84320 0 0 $X=56390 $Y=84080
X240 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 100640 0 0 $X=57770 $Y=100400
X241 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=61640 95200 1 0 $X=61450 $Y=92240
X242 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=62100 116960 0 0 $X=61910 $Y=116720
X243 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=70840 84320 1 0 $X=70650 $Y=81360
X244 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71300 116960 1 0 $X=71110 $Y=114000
X245 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 95200 1 0 $X=72030 $Y=92240
X246 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=81420 89760 0 0 $X=81230 $Y=89520
X247 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=85560 122400 0 0 $X=85370 $Y=122160
X248 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=101200 84320 0 0 $X=101010 $Y=84080
X249 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=111320 100640 0 0 $X=111130 $Y=100400
X250 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=112240 89760 1 0 $X=112050 $Y=86800
X251 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=123740 78880 0 0 $X=123550 $Y=78640
X252 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126960 100640 1 0 $X=126770 $Y=97680
X253 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=127420 95200 1 0 $X=127230 $Y=92240
X254 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=127880 116960 1 0 $X=127690 $Y=114000
X255 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 111520 1 0 $X=132290 $Y=108560
X256 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142140 122400 1 0 $X=141950 $Y=119440
X257 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=151800 100640 0 0 $X=151610 $Y=100400
X258 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 122400 1 0 $X=156210 $Y=119440
X259 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=160540 111520 1 0 $X=160350 $Y=108560
X260 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=161460 116960 0 0 $X=161270 $Y=116720
X261 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 100640 1 0 $X=165410 $Y=97680
X262 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=168820 100640 0 0 $X=168630 $Y=100400
X263 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 95200 1 0 $X=170010 $Y=92240
X264 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=173880 106080 1 0 $X=173690 $Y=103120
X265 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 95200 0 0 $X=174150 $Y=94960
X266 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178020 116960 0 0 $X=177830 $Y=116720
X267 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178940 122400 1 0 $X=178750 $Y=119440
X268 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184000 116960 0 0 $X=183810 $Y=116720
X269 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 106080 1 0 $X=184270 $Y=103120
X270 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 111520 1 0 $X=184270 $Y=108560
X271 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 122400 1 0 $X=184270 $Y=119440
X272 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=195500 100640 1 0 $X=195310 $Y=97680
X273 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=195960 95200 1 0 $X=195770 $Y=92240
X274 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=197340 106080 0 0 $X=197150 $Y=105840
X275 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=199640 106080 1 0 $X=199450 $Y=103120
X276 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 84320 1 0 $X=212330 $Y=81360
X277 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 106080 1 0 $X=212330 $Y=103120
X278 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 95200 1 0 $X=216470 $Y=92240
X279 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=223100 78880 0 0 $X=222910 $Y=78640
X280 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 95200 0 0 $X=226130 $Y=94960
X281 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=228620 106080 1 0 $X=228430 $Y=103120
X282 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 89760 0 0 $X=230270 $Y=89520
X283 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240580 95200 1 0 $X=240390 $Y=92240
X284 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=247480 100640 1 0 $X=247290 $Y=97680
X285 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=252540 100640 0 0 $X=252350 $Y=100400
X286 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258060 100640 1 0 $X=257870 $Y=97680
X287 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281060 100640 0 0 $X=280870 $Y=100400
X288 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=283360 95200 1 0 $X=283170 $Y=92240
X289 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286120 122400 1 0 $X=285930 $Y=119440
X290 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=288420 100640 1 0 $X=288230 $Y=97680
X291 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=291640 111520 0 0 $X=291450 $Y=111280
X292 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=292100 116960 0 0 $X=291910 $Y=116720
X293 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=295320 89760 1 0 $X=295130 $Y=86800
X294 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 100640 1 0 $X=296510 $Y=97680
X295 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=307280 122400 1 0 $X=307090 $Y=119440
X296 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 106080 1 0 $X=310310 $Y=103120
X297 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 111520 1 0 $X=310310 $Y=108560
X298 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=319700 116960 0 0 $X=319510 $Y=116720
X299 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=320160 89760 0 0 $X=319970 $Y=89520
X300 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 106080 1 0 $X=324570 $Y=103120
X301 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 100640 1 0 $X=328710 $Y=97680
X302 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 106080 1 0 $X=328710 $Y=103120
X303 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344080 106080 1 0 $X=343890 $Y=103120
X304 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344540 122400 1 0 $X=344350 $Y=119440
X305 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 84320 1 0 $X=344810 $Y=81360
X306 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 89760 1 0 $X=345270 $Y=86800
X307 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 84320 0 0 $X=6710 $Y=84080
X308 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 89760 1 0 $X=6710 $Y=86800
X309 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 95200 0 0 $X=6710 $Y=94960
X310 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=11040 122400 1 0 $X=10850 $Y=119440
X311 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=18400 78880 0 0 $X=18210 $Y=78640
X312 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=24840 84320 0 0 $X=24650 $Y=84080
X313 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=39100 89760 0 0 $X=38910 $Y=89520
X314 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40480 84320 1 0 $X=40290 $Y=81360
X315 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=52440 116960 1 0 $X=52250 $Y=114000
X316 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=59340 100640 1 0 $X=59150 $Y=97680
X317 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=67160 89760 1 0 $X=66970 $Y=86800
X318 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=68540 116960 0 0 $X=68350 $Y=116720
X319 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=70380 89760 0 0 $X=70190 $Y=89520
X320 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81420 84320 1 0 $X=81230 $Y=81360
X321 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82340 111520 0 0 $X=82150 $Y=111280
X322 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82800 95200 1 0 $X=82610 $Y=92240
X323 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=87860 122400 1 0 $X=87670 $Y=119440
X324 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97520 78880 0 0 $X=97330 $Y=78640
X325 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=98440 84320 1 0 $X=98250 $Y=81360
X326 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=98900 122400 0 0 $X=98710 $Y=122160
X327 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=109480 78880 0 0 $X=109290 $Y=78640
X328 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=110860 122400 0 0 $X=110670 $Y=122160
X329 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=111780 95200 1 0 $X=111590 $Y=92240
X330 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=126040 122400 1 0 $X=125850 $Y=119440
X331 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=126500 84320 1 0 $X=126310 $Y=81360
X332 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=135240 122400 0 0 $X=135050 $Y=122160
X333 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=137540 116960 1 0 $X=137350 $Y=114000
X334 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=139840 100640 0 0 $X=139650 $Y=100400
X335 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=165140 111520 0 0 $X=164950 $Y=111280
X336 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=185380 111520 0 0 $X=185190 $Y=111280
X337 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=190900 111520 1 0 $X=190710 $Y=108560
X338 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=208840 116960 1 0 $X=208650 $Y=114000
X339 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=209760 89760 1 0 $X=209570 $Y=86800
X340 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=217120 111520 0 0 $X=216930 $Y=111280
X341 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=225400 100640 1 0 $X=225210 $Y=97680
X342 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=227700 95200 1 0 $X=227510 $Y=92240
X343 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235520 89760 1 0 $X=235330 $Y=86800
X344 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=247020 95200 1 0 $X=246830 $Y=92240
X345 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=251160 106080 0 0 $X=250970 $Y=105840
X346 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=264960 106080 1 0 $X=264770 $Y=103120
X347 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=290720 111520 1 0 $X=290530 $Y=108560
X348 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=290720 116960 1 0 $X=290530 $Y=114000
X349 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=299000 100640 0 0 $X=298810 $Y=100400
X350 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=320620 111520 1 0 $X=320430 $Y=108560
X351 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=321540 100640 1 0 $X=321350 $Y=97680
X352 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=321540 116960 1 0 $X=321350 $Y=114000
X353 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322460 84320 1 0 $X=322270 $Y=81360
X354 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322920 89760 1 0 $X=322730 $Y=86800
X355 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322920 95200 1 0 $X=322730 $Y=92240
X356 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322920 122400 1 0 $X=322730 $Y=119440
X357 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=323840 106080 0 0 $X=323650 $Y=105840
X358 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=325680 111520 0 0 $X=325490 $Y=111280
X359 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=326140 84320 0 0 $X=325950 $Y=84080
X360 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=326140 100640 0 0 $X=325950 $Y=100400
X361 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=327520 122400 0 0 $X=327330 $Y=122160
X362 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=328900 78880 0 0 $X=328710 $Y=78640
X363 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=342700 111520 1 0 $X=342510 $Y=108560
X364 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=343620 95200 1 0 $X=343430 $Y=92240
X365 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=343620 100640 1 0 $X=343430 $Y=97680
X366 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=343620 116960 1 0 $X=343430 $Y=114000
X367 1 2 ICV_2 $T=33580 78880 0 0 $X=33390 $Y=78640
X368 1 2 ICV_2 $T=75900 89760 1 0 $X=75710 $Y=86800
X369 1 2 ICV_2 $T=103960 84320 1 0 $X=103770 $Y=81360
X370 1 2 ICV_2 $T=117760 78880 0 0 $X=117570 $Y=78640
X371 1 2 ICV_2 $T=145820 100640 0 0 $X=145630 $Y=100400
X372 1 2 ICV_2 $T=145820 106080 0 0 $X=145630 $Y=105840
X373 1 2 ICV_2 $T=145820 116960 0 0 $X=145630 $Y=116720
X374 1 2 ICV_2 $T=173880 106080 0 0 $X=173690 $Y=105840
X375 1 2 ICV_2 $T=188140 116960 1 0 $X=187950 $Y=114000
X376 1 2 ICV_2 $T=216200 106080 1 0 $X=216010 $Y=103120
X377 1 2 ICV_2 $T=216200 111520 1 0 $X=216010 $Y=108560
X378 1 2 ICV_2 $T=286120 100640 0 0 $X=285930 $Y=100400
X379 1 2 ICV_2 $T=286120 116960 0 0 $X=285930 $Y=116720
X380 1 2 ICV_2 $T=314180 89760 0 0 $X=313990 $Y=89520
X381 1 2 ICV_2 $T=328440 84320 1 0 $X=328250 $Y=81360
X382 1 2 ICV_2 $T=342240 78880 0 0 $X=342050 $Y=78640
X383 1 2 ICV_2 $T=342240 84320 0 0 $X=342050 $Y=84080
X384 1 2 ICV_2 $T=342240 89760 0 0 $X=342050 $Y=89520
X385 1 2 ICV_2 $T=342240 95200 0 0 $X=342050 $Y=94960
X386 1 2 ICV_2 $T=342240 100640 0 0 $X=342050 $Y=100400
X387 1 2 ICV_2 $T=342240 106080 0 0 $X=342050 $Y=105840
X388 1 2 ICV_2 $T=342240 111520 0 0 $X=342050 $Y=111280
X389 1 2 ICV_2 $T=342240 116960 0 0 $X=342050 $Y=116720
X390 1 2 ICV_2 $T=342240 122400 0 0 $X=342050 $Y=122160
X391 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 89760 0 0 $X=6710 $Y=89520
X392 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=28060 100640 0 0 $X=27870 $Y=100400
X393 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=28520 122400 0 0 $X=28330 $Y=122160
X394 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 84320 1 0 $X=45810 $Y=81360
X395 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46920 122400 0 0 $X=46730 $Y=122160
X396 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=55200 122400 0 0 $X=55010 $Y=122160
X397 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=57960 116960 1 0 $X=57770 $Y=114000
X398 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59800 122400 0 0 $X=59610 $Y=122160
X399 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=64860 100640 1 0 $X=64670 $Y=97680
X400 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73140 100640 0 0 $X=72950 $Y=100400
X401 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=74060 116960 0 0 $X=73870 $Y=116720
X402 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 100640 1 0 $X=76170 $Y=97680
X403 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=85560 78880 0 0 $X=85370 $Y=78640
X404 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=86020 106080 1 0 $X=85830 $Y=103120
X405 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87400 84320 0 0 $X=87210 $Y=84080
X406 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87860 111520 0 0 $X=87670 $Y=111280
X407 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=92000 89760 1 0 $X=91810 $Y=86800
X408 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=101660 111520 1 0 $X=101470 $Y=108560
X409 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 116960 0 0 $X=104230 $Y=116720
X410 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=106720 100640 0 0 $X=106530 $Y=100400
X411 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=112700 106080 1 0 $X=112510 $Y=103120
X412 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115460 100640 1 0 $X=115270 $Y=97680
X413 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=117300 89760 1 0 $X=117110 $Y=86800
X414 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=121440 84320 0 0 $X=121250 $Y=84080
X415 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=130180 111520 1 0 $X=129990 $Y=108560
X416 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=137540 84320 1 0 $X=137350 $Y=81360
X417 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=148580 84320 0 0 $X=148390 $Y=84080
X418 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=151340 89760 0 0 $X=151150 $Y=89520
X419 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=154100 89760 1 0 $X=153910 $Y=86800
X420 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 116960 1 0 $X=160350 $Y=114000
X421 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 78880 0 0 $X=171850 $Y=78640
X422 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=187680 95200 0 0 $X=187490 $Y=94960
X423 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=192740 95200 1 0 $X=192550 $Y=92240
X424 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=195040 122400 1 0 $X=194850 $Y=119440
X425 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=195960 111520 0 0 $X=195770 $Y=111280
X426 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=199640 122400 0 0 $X=199450 $Y=122160
X427 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=204700 89760 0 0 $X=204510 $Y=89520
X428 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=206080 106080 1 0 $X=205890 $Y=103120
X429 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=207460 78880 0 0 $X=207270 $Y=78640
X430 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 116960 1 0 $X=214170 $Y=114000
X431 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216200 116960 0 0 $X=216010 $Y=116720
X432 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=222640 111520 0 0 $X=222450 $Y=111280
X433 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=227700 84320 0 0 $X=227510 $Y=84080
X434 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230000 84320 1 0 $X=229810 $Y=81360
X435 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230000 122400 1 0 $X=229810 $Y=119440
X436 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=234600 95200 0 0 $X=234410 $Y=94960
X437 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=243800 111520 0 0 $X=243610 $Y=111280
X438 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=246100 116960 0 0 $X=245910 $Y=116720
X439 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=250240 89760 0 0 $X=250050 $Y=89520
X440 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=253920 84320 1 0 $X=253730 $Y=81360
X441 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=261280 84320 1 0 $X=261090 $Y=81360
X442 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=270480 84320 0 0 $X=270290 $Y=84080
X443 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=270480 106080 1 0 $X=270290 $Y=103120
X444 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=281980 95200 0 0 $X=281790 $Y=94960
X445 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=296240 111520 1 0 $X=296050 $Y=108560
X446 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=296240 116960 1 0 $X=296050 $Y=114000
X447 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=296240 122400 1 0 $X=296050 $Y=119440
X448 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=297620 78880 0 0 $X=297430 $Y=78640
X449 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=299460 89760 0 0 $X=299270 $Y=89520
X450 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=304520 100640 0 0 $X=304330 $Y=100400
X451 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=304980 89760 1 0 $X=304790 $Y=86800
X452 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=310040 84320 0 0 $X=309850 $Y=84080
X453 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=314640 122400 0 0 $X=314450 $Y=122160
X454 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=315100 100640 1 0 $X=314910 $Y=97680
X455 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 111520 1 0 $X=325950 $Y=108560
X456 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=331200 111520 0 0 $X=331010 $Y=111280
X457 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=331660 100640 0 0 $X=331470 $Y=100400
X458 1 12 sky130_fd_sc_hd__diode_2 $T=7820 122400 1 0 $X=7630 $Y=119440
X459 1 12 sky130_fd_sc_hd__diode_2 $T=12420 84320 0 0 $X=12230 $Y=84080
X460 1 17 sky130_fd_sc_hd__diode_2 $T=19320 116960 0 0 $X=19130 $Y=116720
X461 1 24 sky130_fd_sc_hd__diode_2 $T=22540 95200 1 0 $X=22350 $Y=92240
X462 1 415 sky130_fd_sc_hd__diode_2 $T=23920 78880 0 0 $X=23730 $Y=78640
X463 1 413 sky130_fd_sc_hd__diode_2 $T=34960 106080 0 0 $X=34770 $Y=105840
X464 1 39 sky130_fd_sc_hd__diode_2 $T=41400 100640 0 0 $X=41210 $Y=100400
X465 1 42 sky130_fd_sc_hd__diode_2 $T=43700 122400 0 0 $X=43510 $Y=122160
X466 1 430 sky130_fd_sc_hd__diode_2 $T=49220 95200 1 0 $X=49030 $Y=92240
X467 1 441 sky130_fd_sc_hd__diode_2 $T=49220 116960 1 0 $X=49030 $Y=114000
X468 1 45 sky130_fd_sc_hd__diode_2 $T=49220 122400 0 0 $X=49030 $Y=122160
X469 1 12 sky130_fd_sc_hd__diode_2 $T=49680 89760 0 0 $X=49490 $Y=89520
X470 1 439 sky130_fd_sc_hd__diode_2 $T=67620 106080 0 0 $X=67430 $Y=105840
X471 1 60 sky130_fd_sc_hd__diode_2 $T=68080 78880 0 0 $X=67890 $Y=78640
X472 1 68 sky130_fd_sc_hd__diode_2 $T=77280 122400 0 0 $X=77090 $Y=122160
X473 1 72 sky130_fd_sc_hd__diode_2 $T=82340 78880 0 0 $X=82150 $Y=78640
X474 1 466 sky130_fd_sc_hd__diode_2 $T=92000 106080 1 0 $X=91810 $Y=103120
X475 1 474 sky130_fd_sc_hd__diode_2 $T=92000 116960 1 0 $X=91810 $Y=114000
X476 1 75 sky130_fd_sc_hd__diode_2 $T=92460 111520 0 0 $X=92270 $Y=111280
X477 1 80 sky130_fd_sc_hd__diode_2 $T=95220 84320 0 0 $X=95030 $Y=84080
X478 1 83 sky130_fd_sc_hd__diode_2 $T=95220 89760 0 0 $X=95030 $Y=89520
X479 1 458 sky130_fd_sc_hd__diode_2 $T=99360 89760 0 0 $X=99170 $Y=89520
X480 1 85 sky130_fd_sc_hd__diode_2 $T=103500 78880 0 0 $X=103310 $Y=78640
X481 1 483 sky130_fd_sc_hd__diode_2 $T=106720 116960 1 0 $X=106530 $Y=114000
X482 1 487 sky130_fd_sc_hd__diode_2 $T=113620 106080 0 0 $X=113430 $Y=105840
X483 1 472 sky130_fd_sc_hd__diode_2 $T=119140 95200 0 0 $X=118950 $Y=94960
X484 1 97 sky130_fd_sc_hd__diode_2 $T=120980 100640 1 0 $X=120790 $Y=97680
X485 1 112 sky130_fd_sc_hd__diode_2 $T=133860 100640 0 0 $X=133670 $Y=100400
X486 1 502 sky130_fd_sc_hd__diode_2 $T=134320 89760 0 0 $X=134130 $Y=89520
X487 1 115 sky130_fd_sc_hd__diode_2 $T=136160 78880 0 0 $X=135970 $Y=78640
X488 1 499 sky130_fd_sc_hd__diode_2 $T=138000 89760 1 0 $X=137810 $Y=86800
X489 1 504 sky130_fd_sc_hd__diode_2 $T=141680 84320 0 0 $X=141490 $Y=84080
X490 1 491 sky130_fd_sc_hd__diode_2 $T=147200 111520 0 0 $X=147010 $Y=111280
X491 1 503 sky130_fd_sc_hd__diode_2 $T=152260 106080 0 0 $X=152070 $Y=105840
X492 1 507 sky130_fd_sc_hd__diode_2 $T=153640 89760 0 0 $X=153450 $Y=89520
X493 1 130 sky130_fd_sc_hd__diode_2 $T=154100 84320 0 0 $X=153910 $Y=84080
X494 1 134 sky130_fd_sc_hd__diode_2 $T=155480 100640 0 0 $X=155290 $Y=100400
X495 1 135 sky130_fd_sc_hd__diode_2 $T=158700 122400 0 0 $X=158510 $Y=122160
X496 1 397 sky130_fd_sc_hd__diode_2 $T=171120 89760 1 0 $X=170930 $Y=86800
X497 1 519 sky130_fd_sc_hd__diode_2 $T=179400 84320 0 0 $X=179210 $Y=84080
X498 1 156 sky130_fd_sc_hd__diode_2 $T=181700 89760 0 0 $X=181510 $Y=89520
X499 1 145 sky130_fd_sc_hd__diode_2 $T=189520 84320 1 0 $X=189330 $Y=81360
X500 1 157 sky130_fd_sc_hd__diode_2 $T=189980 95200 0 0 $X=189790 $Y=94960
X501 1 12 sky130_fd_sc_hd__diode_2 $T=206540 106080 0 0 $X=206350 $Y=105840
X502 1 12 sky130_fd_sc_hd__diode_2 $T=207000 89760 0 0 $X=206810 $Y=89520
X503 1 177 sky130_fd_sc_hd__diode_2 $T=210680 116960 0 0 $X=210490 $Y=116720
X504 1 182 sky130_fd_sc_hd__diode_2 $T=211600 122400 0 0 $X=211410 $Y=122160
X505 1 185 sky130_fd_sc_hd__diode_2 $T=217120 100640 0 0 $X=216930 $Y=100400
X506 1 185 sky130_fd_sc_hd__diode_2 $T=225860 122400 0 0 $X=225670 $Y=122160
X507 1 12 sky130_fd_sc_hd__diode_2 $T=231380 106080 0 0 $X=231190 $Y=105840
X508 1 207 sky130_fd_sc_hd__diode_2 $T=236900 95200 0 0 $X=236710 $Y=94960
X509 1 543 sky130_fd_sc_hd__diode_2 $T=244260 89760 0 0 $X=244070 $Y=89520
X510 1 213 sky130_fd_sc_hd__diode_2 $T=245640 84320 1 0 $X=245450 $Y=81360
X511 1 217 sky130_fd_sc_hd__diode_2 $T=248400 116960 0 0 $X=248210 $Y=116720
X512 1 538 sky130_fd_sc_hd__diode_2 $T=253920 111520 0 0 $X=253730 $Y=111280
X513 1 222 sky130_fd_sc_hd__diode_2 $T=264500 78880 0 0 $X=264310 $Y=78640
X514 1 227 sky130_fd_sc_hd__diode_2 $T=264500 84320 0 0 $X=264310 $Y=84080
X515 1 230 sky130_fd_sc_hd__diode_2 $T=268180 84320 1 0 $X=267990 $Y=81360
X516 1 556 sky130_fd_sc_hd__diode_2 $T=268180 89760 0 0 $X=267990 $Y=89520
X517 1 234 sky130_fd_sc_hd__diode_2 $T=272320 122400 0 0 $X=272130 $Y=122160
X518 1 561 sky130_fd_sc_hd__diode_2 $T=272780 111520 0 0 $X=272590 $Y=111280
X519 1 169 sky130_fd_sc_hd__diode_2 $T=273700 116960 1 0 $X=273510 $Y=114000
X520 1 235 sky130_fd_sc_hd__diode_2 $T=276000 84320 0 0 $X=275810 $Y=84080
X521 1 233 sky130_fd_sc_hd__diode_2 $T=277380 95200 1 0 $X=277190 $Y=92240
X522 1 235 sky130_fd_sc_hd__diode_2 $T=279220 84320 1 0 $X=279030 $Y=81360
X523 1 244 sky130_fd_sc_hd__diode_2 $T=292560 78880 0 0 $X=292370 $Y=78640
X524 1 559 sky130_fd_sc_hd__diode_2 $T=292560 89760 0 0 $X=292370 $Y=89520
X525 1 571 sky130_fd_sc_hd__diode_2 $T=293020 100640 0 0 $X=292830 $Y=100400
X526 1 252 sky130_fd_sc_hd__diode_2 $T=300840 116960 0 0 $X=300650 $Y=116720
X527 1 242 sky130_fd_sc_hd__diode_2 $T=301760 89760 0 0 $X=301570 $Y=89520
X528 1 252 sky130_fd_sc_hd__diode_2 $T=301760 106080 1 0 $X=301570 $Y=103120
X529 1 544 sky130_fd_sc_hd__diode_2 $T=304980 84320 0 0 $X=304790 $Y=84080
X530 1 577 sky130_fd_sc_hd__diode_2 $T=308200 116960 1 0 $X=308010 $Y=114000
X531 1 258 sky130_fd_sc_hd__diode_2 $T=310040 89760 1 0 $X=309850 $Y=86800
X532 1 582 sky130_fd_sc_hd__diode_2 $T=310500 84320 1 0 $X=310310 $Y=81360
X533 1 586 sky130_fd_sc_hd__diode_2 $T=331200 95200 1 0 $X=331010 $Y=92240
X534 1 11 sky130_fd_sc_hd__diode_2 $T=333040 89760 1 0 $X=332850 $Y=86800
X535 1 2 420 ICV_4 $T=26220 111520 1 0 $X=26030 $Y=108560
X536 1 2 29 ICV_4 $T=30360 84320 0 0 $X=30170 $Y=84080
X537 1 2 12 ICV_4 $T=30820 78880 0 0 $X=30630 $Y=78640
X538 1 2 30 ICV_4 $T=30820 122400 0 0 $X=30630 $Y=122160
X539 1 2 433 ICV_4 $T=46460 111520 0 0 $X=46270 $Y=111280
X540 1 2 12 ICV_4 $T=48300 78880 0 0 $X=48110 $Y=78640
X541 1 2 438 ICV_4 $T=51060 106080 0 0 $X=50870 $Y=105840
X542 1 2 438 ICV_4 $T=56580 95200 0 0 $X=56390 $Y=94960
X543 1 2 50 ICV_4 $T=58420 106080 0 0 $X=58230 $Y=105840
X544 1 2 429 ICV_4 $T=58880 89760 0 0 $X=58690 $Y=89520
X545 1 2 58 ICV_4 $T=73140 106080 1 0 $X=72950 $Y=103120
X546 1 2 456 ICV_4 $T=76360 111520 0 0 $X=76170 $Y=111280
X547 1 2 445 ICV_4 $T=76820 106080 0 0 $X=76630 $Y=105840
X548 1 2 466 ICV_4 $T=83720 100640 1 0 $X=83530 $Y=97680
X549 1 2 51 ICV_4 $T=86940 106080 0 0 $X=86750 $Y=105840
X550 1 2 472 ICV_4 $T=91540 100640 1 0 $X=91350 $Y=97680
X551 1 2 468 ICV_4 $T=96140 106080 0 0 $X=95950 $Y=105840
X552 1 2 475 ICV_4 $T=96140 111520 1 0 $X=95950 $Y=108560
X553 1 2 479 ICV_4 $T=101200 95200 1 0 $X=101010 $Y=92240
X554 1 2 476 ICV_4 $T=101200 106080 1 0 $X=101010 $Y=103120
X555 1 2 84 ICV_4 $T=105340 106080 1 0 $X=105150 $Y=103120
X556 1 2 77 ICV_4 $T=106720 116960 0 0 $X=106530 $Y=116720
X557 1 2 94 ICV_4 $T=113620 111520 1 0 $X=113430 $Y=108560
X558 1 2 93 ICV_4 $T=115000 84320 0 0 $X=114810 $Y=84080
X559 1 2 483 ICV_4 $T=115000 111520 0 0 $X=114810 $Y=111280
X560 1 2 486 ICV_4 $T=115000 116960 0 0 $X=114810 $Y=116720
X561 1 2 462 ICV_4 $T=119140 106080 0 0 $X=118950 $Y=105840
X562 1 2 115 ICV_4 $T=141220 89760 0 0 $X=141030 $Y=89520
X563 1 2 502 ICV_4 $T=141220 95200 0 0 $X=141030 $Y=94960
X564 1 2 501 ICV_4 $T=143060 78880 0 0 $X=142870 $Y=78640
X565 1 2 500 ICV_4 $T=147200 100640 1 0 $X=147010 $Y=97680
X566 1 2 504 ICV_4 $T=149960 89760 1 0 $X=149770 $Y=86800
X567 1 2 112 ICV_4 $T=151340 95200 1 0 $X=151150 $Y=92240
X568 1 2 115 ICV_4 $T=151800 95200 0 0 $X=151610 $Y=94960
X569 1 2 107 ICV_4 $T=152260 84320 1 0 $X=152070 $Y=81360
X570 1 2 122 ICV_4 $T=155940 78880 0 0 $X=155750 $Y=78640
X571 1 2 131 ICV_4 $T=156860 95200 0 0 $X=156670 $Y=94960
X572 1 2 504 ICV_4 $T=157320 84320 1 0 $X=157130 $Y=81360
X573 1 2 115 ICV_4 $T=160540 89760 0 0 $X=160350 $Y=89520
X574 1 2 464 ICV_4 $T=166520 84320 1 0 $X=166330 $Y=81360
X575 1 2 498 ICV_4 $T=177100 84320 1 0 $X=176910 $Y=81360
X576 1 2 109 ICV_4 $T=186300 84320 0 0 $X=186110 $Y=84080
X577 1 2 122 ICV_4 $T=193200 84320 0 0 $X=193010 $Y=84080
X578 1 2 389 ICV_4 $T=193200 89760 1 0 $X=193010 $Y=86800
X579 1 2 165 ICV_4 $T=193660 116960 0 0 $X=193470 $Y=116720
X580 1 2 521 ICV_4 $T=196880 95200 0 0 $X=196690 $Y=94960
X581 1 2 6 ICV_4 $T=199640 84320 1 0 $X=199450 $Y=81360
X582 1 2 7 ICV_4 $T=199640 95200 1 0 $X=199450 $Y=92240
X583 1 2 523 ICV_4 $T=200100 89760 1 0 $X=199910 $Y=86800
X584 1 2 167 ICV_4 $T=203320 106080 0 0 $X=203130 $Y=105840
X585 1 2 176 ICV_4 $T=206540 84320 1 0 $X=206350 $Y=81360
X586 1 2 158 ICV_4 $T=208380 122400 0 0 $X=208190 $Y=122160
X587 1 2 184 ICV_4 $T=221720 116960 0 0 $X=221530 $Y=116720
X588 1 2 187 ICV_4 $T=224480 122400 1 0 $X=224290 $Y=119440
X589 1 2 191 ICV_4 $T=227240 111520 0 0 $X=227050 $Y=111280
X590 1 2 537 ICV_4 $T=230920 89760 1 0 $X=230730 $Y=86800
X591 1 2 540 ICV_4 $T=233220 106080 1 0 $X=233030 $Y=103120
X592 1 2 191 ICV_4 $T=239660 111520 0 0 $X=239470 $Y=111280
X593 1 2 209 ICV_4 $T=241500 84320 1 0 $X=241310 $Y=81360
X594 1 2 214 ICV_4 $T=245640 89760 1 0 $X=245450 $Y=86800
X595 1 2 216 ICV_4 $T=251620 78880 0 0 $X=251430 $Y=78640
X596 1 2 213 ICV_4 $T=260360 89760 1 0 $X=260170 $Y=86800
X597 1 2 546 ICV_4 $T=262660 95200 1 0 $X=262470 $Y=92240
X598 1 2 557 ICV_4 $T=265420 89760 1 0 $X=265230 $Y=86800
X599 1 2 227 ICV_4 $T=270480 78880 0 0 $X=270290 $Y=78640
X600 1 2 548 ICV_4 $T=272780 84320 0 0 $X=272590 $Y=84080
X601 1 2 221 ICV_4 $T=276000 84320 1 0 $X=275810 $Y=81360
X602 1 2 226 ICV_4 $T=281520 122400 0 0 $X=281330 $Y=122160
X603 1 2 235 ICV_4 $T=282900 84320 0 0 $X=282710 $Y=84080
X604 1 2 233 ICV_4 $T=289340 95200 1 0 $X=289150 $Y=92240
X605 1 2 258 ICV_4 $T=306820 89760 1 0 $X=306630 $Y=86800
X606 1 2 259 ICV_4 $T=307740 84320 1 0 $X=307550 $Y=81360
X607 1 2 266 ICV_4 $T=316940 89760 1 0 $X=316750 $Y=86800
X608 1 2 587 ICV_4 $T=329820 89760 1 0 $X=329630 $Y=86800
X609 1 2 272 ICV_4 $T=329820 116960 1 0 $X=329630 $Y=114000
X610 1 2 12 ICV_4 $T=339480 89760 0 0 $X=339290 $Y=89520
X611 1 2 11 ICV_4 $T=339480 116960 0 0 $X=339290 $Y=116720
X612 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 100640 1 0 $X=16370 $Y=97680
X613 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 122400 1 0 $X=16370 $Y=119440
X614 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=18400 100640 0 0 $X=18210 $Y=100400
X615 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=28980 116960 0 0 $X=28790 $Y=116720
X616 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=40480 106080 1 0 $X=40290 $Y=103120
X617 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 89760 1 0 $X=72490 $Y=86800
X618 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 122400 1 0 $X=72490 $Y=119440
X619 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 111520 0 0 $X=72950 $Y=111280
X620 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=75900 89760 0 0 $X=75710 $Y=89520
X621 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=79120 78880 0 0 $X=78930 $Y=78640
X622 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=81880 89760 1 0 $X=81690 $Y=86800
X623 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=89700 111520 1 0 $X=89510 $Y=108560
X624 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=100740 116960 1 0 $X=100550 $Y=114000
X625 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=108100 89760 1 0 $X=107910 $Y=86800
X626 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 78880 0 0 $X=114810 $Y=78640
X627 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=118220 122400 0 0 $X=118030 $Y=122160
X628 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=126040 84320 0 0 $X=125850 $Y=84080
X629 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 106080 1 0 $X=132290 $Y=103120
X630 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=140760 122400 0 0 $X=140570 $Y=122160
X631 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=142600 106080 0 0 $X=142410 $Y=105840
X632 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=151800 116960 0 0 $X=151610 $Y=116720
X633 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=170660 111520 0 0 $X=170470 $Y=111280
X634 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=171120 106080 0 0 $X=170930 $Y=105840
X635 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=177100 111520 1 0 $X=176910 $Y=108560
X636 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185840 122400 0 0 $X=185650 $Y=122160
X637 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=186760 106080 0 0 $X=186570 $Y=105840
X638 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=190900 122400 1 0 $X=190710 $Y=119440
X639 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 106080 0 0 $X=226590 $Y=105840
X640 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=227700 89760 1 0 $X=227510 $Y=86800
X641 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=228620 111520 1 0 $X=228430 $Y=108560
X642 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=233220 95200 1 0 $X=233030 $Y=92240
X643 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=235980 100640 1 0 $X=235790 $Y=97680
X644 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241040 89760 1 0 $X=240850 $Y=86800
X645 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241500 122400 1 0 $X=241310 $Y=119440
X646 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 122400 1 0 $X=244530 $Y=119440
X647 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=248400 111520 0 0 $X=248210 $Y=111280
X648 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=255760 106080 1 0 $X=255570 $Y=103120
X649 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=258520 95200 0 0 $X=258330 $Y=94960
X650 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=270020 111520 0 0 $X=269830 $Y=111280
X651 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=272780 111520 1 0 $X=272590 $Y=108560
X652 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=279220 122400 1 0 $X=279030 $Y=119440
X653 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=282900 106080 0 0 $X=282710 $Y=105840
X654 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=284280 100640 1 0 $X=284090 $Y=97680
X655 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297160 95200 1 0 $X=296970 $Y=92240
X656 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=298080 84320 0 0 $X=297890 $Y=84080
X657 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=298080 122400 0 0 $X=297890 $Y=122160
X658 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=310960 95200 0 0 $X=310770 $Y=94960
X659 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 95200 0 0 $X=314450 $Y=94960
X660 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=328900 111520 1 0 $X=328710 $Y=108560
X661 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=329360 106080 0 0 $X=329170 $Y=105840
X662 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331660 84320 0 0 $X=331470 $Y=84080
X663 1 2 25 ICV_5 $T=26220 89760 1 0 $X=26030 $Y=86800
X664 1 2 424 ICV_5 $T=28060 89760 0 0 $X=27870 $Y=89520
X665 1 2 422 ICV_5 $T=29900 111520 0 0 $X=29710 $Y=111280
X666 1 2 423 ICV_5 $T=40020 111520 0 0 $X=39830 $Y=111280
X667 1 2 419 ICV_5 $T=41400 95200 0 0 $X=41210 $Y=94960
X668 1 2 432 ICV_5 $T=43700 116960 1 0 $X=43510 $Y=114000
X669 1 2 36 ICV_5 $T=54280 111520 0 0 $X=54090 $Y=111280
X670 1 2 462 ICV_5 $T=84640 111520 1 0 $X=84450 $Y=108560
X671 1 2 98 ICV_5 $T=115920 84320 1 0 $X=115730 $Y=81360
X672 1 2 105 ICV_5 $T=128800 122400 0 0 $X=128610 $Y=122160
X673 1 2 126 ICV_5 $T=150880 122400 1 0 $X=150690 $Y=119440
X674 1 2 168 ICV_5 $T=208380 95200 0 0 $X=208190 $Y=94960
X675 1 2 198 ICV_5 $T=232300 84320 1 0 $X=232110 $Y=81360
X676 1 2 277 ICV_5 $T=338100 78880 0 0 $X=337910 $Y=78640
X677 1 2 281 ICV_5 $T=338100 122400 0 0 $X=337910 $Y=122160
X678 1 2 278 ICV_5 $T=338560 84320 0 0 $X=338370 $Y=84080
X679 1 2 409 ICV_6 $T=14260 84320 1 0 $X=14070 $Y=81360
X680 1 2 411 ICV_6 $T=21160 111520 1 0 $X=20970 $Y=108560
X681 1 2 412 ICV_6 $T=21160 116960 1 0 $X=20970 $Y=114000
X682 1 2 416 ICV_6 $T=23920 106080 1 0 $X=23730 $Y=103120
X683 1 2 41 ICV_6 $T=43240 100640 1 0 $X=43050 $Y=97680
X684 1 2 431 ICV_6 $T=43240 106080 1 0 $X=43050 $Y=103120
X685 1 2 41 ICV_6 $T=49220 111520 1 0 $X=49030 $Y=108560
X686 1 2 429 ICV_6 $T=54280 111520 1 0 $X=54090 $Y=108560
X687 1 2 70 ICV_6 $T=80040 84320 0 0 $X=79850 $Y=84080
X688 1 2 84 ICV_6 $T=98440 122400 1 0 $X=98250 $Y=119440
X689 1 2 459 ICV_6 $T=98900 89760 1 0 $X=98710 $Y=86800
X690 1 2 89 ICV_6 $T=110860 84320 1 0 $X=110670 $Y=81360
X691 1 2 484 ICV_6 $T=115920 116960 1 0 $X=115730 $Y=114000
X692 1 2 495 ICV_6 $T=127420 106080 1 0 $X=127230 $Y=103120
X693 1 2 105 ICV_6 $T=139840 116960 0 0 $X=139650 $Y=116720
X694 1 2 121 ICV_6 $T=146280 122400 1 0 $X=146090 $Y=119440
X695 1 2 130 ICV_6 $T=165600 89760 0 0 $X=165410 $Y=89520
X696 1 2 145 ICV_6 $T=166520 89760 1 0 $X=166330 $Y=86800
X697 1 2 147 ICV_6 $T=169280 116960 0 0 $X=169090 $Y=116720
X698 1 2 517 ICV_6 $T=174340 95200 1 0 $X=174150 $Y=92240
X699 1 2 87 ICV_6 $T=183540 95200 1 0 $X=183350 $Y=92240
X700 1 2 42 ICV_6 $T=188600 116960 0 0 $X=188410 $Y=116720
X701 1 2 156 ICV_6 $T=194580 89760 0 0 $X=194390 $Y=89520
X702 1 2 36 ICV_6 $T=198720 111520 1 0 $X=198530 $Y=108560
X703 1 2 181 ICV_6 $T=212520 100640 0 0 $X=212330 $Y=100400
X704 1 2 539 ICV_6 $T=231840 111520 1 0 $X=231650 $Y=108560
X705 1 2 199 ICV_6 $T=236440 84320 0 0 $X=236250 $Y=84080
X706 1 2 536 ICV_6 $T=236900 116960 1 0 $X=236710 $Y=114000
X707 1 2 537 ICV_6 $T=238740 100640 1 0 $X=238550 $Y=97680
X708 1 2 552 ICV_6 $T=264500 122400 1 0 $X=264310 $Y=119440
X709 1 2 218 ICV_6 $T=264960 116960 1 0 $X=264770 $Y=114000
X710 1 2 559 ICV_6 $T=266800 100640 1 0 $X=266610 $Y=97680
X711 1 2 228 ICV_6 $T=267720 95200 1 0 $X=267530 $Y=92240
X712 1 2 562 ICV_6 $T=275540 111520 1 0 $X=275350 $Y=108560
X713 1 2 191 ICV_6 $T=279220 111520 0 0 $X=279030 $Y=111280
X714 1 2 546 ICV_6 $T=294860 106080 1 0 $X=294670 $Y=103120
X715 1 2 198 ICV_6 $T=295320 84320 1 0 $X=295130 $Y=81360
X716 1 2 275 ICV_6 $T=336720 95200 0 0 $X=336530 $Y=94960
X717 1 2 276 ICV_6 $T=336720 111520 0 0 $X=336530 $Y=111280
X718 1 2 271 ICV_6 $T=337180 100640 0 0 $X=336990 $Y=100400
X719 1 11 12 ICV_7 $T=7820 100640 1 0 $X=7630 $Y=97680
X720 1 11 14 ICV_7 $T=7820 106080 1 0 $X=7630 $Y=103120
X721 1 12 15 ICV_7 $T=7820 111520 1 0 $X=7630 $Y=108560
X722 1 11 16 ICV_7 $T=7820 116960 1 0 $X=7630 $Y=114000
X723 1 17 12 ICV_7 $T=9200 89760 0 0 $X=9010 $Y=89520
X724 1 407 408 ICV_7 $T=12880 89760 1 0 $X=12690 $Y=86800
X725 1 17 414 ICV_7 $T=21160 84320 1 0 $X=20970 $Y=81360
X726 1 413 25 ICV_7 $T=21620 100640 0 0 $X=21430 $Y=100400
X727 1 24 419 ICV_7 $T=24380 89760 0 0 $X=24190 $Y=89520
X728 1 418 421 ICV_7 $T=25300 100640 0 0 $X=25110 $Y=100400
X729 1 24 25 ICV_7 $T=26220 111520 0 0 $X=26030 $Y=111280
X730 1 12 417 ICV_7 $T=26220 116960 0 0 $X=26030 $Y=116720
X731 1 422 28 ICV_7 $T=27600 106080 0 0 $X=27410 $Y=105840
X732 1 427 38 ICV_7 $T=35880 84320 0 0 $X=35690 $Y=84080
X733 1 426 426 ICV_7 $T=35880 95200 1 0 $X=35690 $Y=92240
X734 1 35 40 ICV_7 $T=36340 111520 0 0 $X=36150 $Y=111280
X735 1 435 439 ICV_7 $T=45080 95200 0 0 $X=44890 $Y=94960
X736 1 44 46 ICV_7 $T=48760 95200 0 0 $X=48570 $Y=94960
X737 1 46 439 ICV_7 $T=53360 89760 1 0 $X=53170 $Y=86800
X738 1 41 442 ICV_7 $T=53820 84320 0 0 $X=53630 $Y=84080
X739 1 438 48 ICV_7 $T=55200 100640 0 0 $X=55010 $Y=100400
X740 1 50 51 ICV_7 $T=57040 122400 0 0 $X=56850 $Y=122160
X741 1 55 53 ICV_7 $T=60720 84320 1 0 $X=60530 $Y=81360
X742 1 439 448 ICV_7 $T=62100 111520 1 0 $X=61910 $Y=108560
X743 1 445 430 ICV_7 $T=63020 100640 0 0 $X=62830 $Y=100400
X744 1 446 445 ICV_7 $T=63940 89760 0 0 $X=63750 $Y=89520
X745 1 447 59 ICV_7 $T=63940 106080 1 0 $X=63750 $Y=103120
X746 1 58 439 ICV_7 $T=63940 106080 0 0 $X=63750 $Y=105840
X747 1 50 62 ICV_7 $T=65780 116960 0 0 $X=65590 $Y=116720
X748 1 449 450 ICV_7 $T=66700 100640 1 0 $X=66510 $Y=97680
X749 1 429 451 ICV_7 $T=67620 89760 0 0 $X=67430 $Y=89520
X750 1 50 66 ICV_7 $T=69920 122400 1 0 $X=69730 $Y=119440
X751 1 57 452 ICV_7 $T=70380 100640 1 0 $X=70190 $Y=97680
X752 1 66 454 ICV_7 $T=70380 111520 0 0 $X=70190 $Y=111280
X753 1 66 445 ICV_7 $T=74980 100640 0 0 $X=74790 $Y=100400
X754 1 12 453 ICV_7 $T=76360 116960 0 0 $X=76170 $Y=116720
X755 1 460 463 ICV_7 $T=78660 89760 0 0 $X=78470 $Y=89520
X756 1 460 464 ICV_7 $T=78660 95200 0 0 $X=78470 $Y=94960
X757 1 461 459 ICV_7 $T=79580 111520 0 0 $X=79390 $Y=111280
X758 1 465 467 ICV_7 $T=82340 95200 0 0 $X=82150 $Y=94960
X759 1 73 61 ICV_7 $T=84640 84320 0 0 $X=84450 $Y=84080
X760 1 459 464 ICV_7 $T=88320 106080 1 0 $X=88130 $Y=103120
X761 1 470 77 ICV_7 $T=91080 122400 0 0 $X=90890 $Y=122160
X762 1 76 78 ICV_7 $T=92460 111520 1 0 $X=92270 $Y=108560
X763 1 64 76 ICV_7 $T=95220 100640 0 0 $X=95030 $Y=100400
X764 1 468 446 ICV_7 $T=96140 95200 0 0 $X=95950 $Y=94960
X765 1 475 478 ICV_7 $T=97980 116960 1 0 $X=97790 $Y=114000
X766 1 477 476 ICV_7 $T=98440 100640 1 0 $X=98250 $Y=97680
X767 1 83 464 ICV_7 $T=98900 100640 0 0 $X=98710 $Y=100400
X768 1 450 476 ICV_7 $T=98900 111520 1 0 $X=98710 $Y=108560
X769 1 475 475 ICV_7 $T=103960 111520 0 0 $X=103770 $Y=111280
X770 1 83 479 ICV_7 $T=105340 89760 1 0 $X=105150 $Y=86800
X771 1 461 476 ICV_7 $T=106260 106080 0 0 $X=106070 $Y=105840
X772 1 475 480 ICV_7 $T=108560 89760 0 0 $X=108370 $Y=89520
X773 1 466 83 ICV_7 $T=108560 100640 0 0 $X=108370 $Y=100400
X774 1 482 94 ICV_7 $T=109940 106080 0 0 $X=109750 $Y=105840
X775 1 96 485 ICV_7 $T=111780 122400 1 0 $X=111590 $Y=119440
X776 1 483 489 ICV_7 $T=112240 89760 0 0 $X=112050 $Y=89520
X777 1 490 95 ICV_7 $T=114540 106080 1 0 $X=114350 $Y=103120
X778 1 99 101 ICV_7 $T=117300 95200 1 0 $X=117110 $Y=92240
X779 1 492 100 ICV_7 $T=117300 100640 1 0 $X=117110 $Y=97680
X780 1 101 465 ICV_7 $T=119140 89760 0 0 $X=118950 $Y=89520
X781 1 467 483 ICV_7 $T=119140 100640 0 0 $X=118950 $Y=100400
X782 1 95 488 ICV_7 $T=119140 111520 0 0 $X=118950 $Y=111280
X783 1 103 483 ICV_7 $T=119600 89760 1 0 $X=119410 $Y=86800
X784 1 479 105 ICV_7 $T=120980 122400 0 0 $X=120790 $Y=122160
X785 1 89 100 ICV_7 $T=123280 84320 0 0 $X=123090 $Y=84080
X786 1 96 103 ICV_7 $T=123740 106080 1 0 $X=123550 $Y=103120
X787 1 494 497 ICV_7 $T=128340 89760 1 0 $X=128150 $Y=86800
X788 1 108 109 ICV_7 $T=129260 84320 0 0 $X=129070 $Y=84080
X789 1 491 499 ICV_7 $T=130180 100640 0 0 $X=129990 $Y=100400
X790 1 498 113 ICV_7 $T=132480 78880 0 0 $X=132290 $Y=78640
X791 1 501 502 ICV_7 $T=132480 95200 0 0 $X=132290 $Y=94960
X792 1 105 94 ICV_7 $T=132480 122400 0 0 $X=132290 $Y=122160
X793 1 499 112 ICV_7 $T=132940 84320 0 0 $X=132750 $Y=84080
X794 1 111 499 ICV_7 $T=133400 100640 1 0 $X=133210 $Y=97680
X795 1 499 501 ICV_7 $T=134320 89760 1 0 $X=134130 $Y=86800
X796 1 111 112 ICV_7 $T=134320 95200 1 0 $X=134130 $Y=92240
X797 1 114 500 ICV_7 $T=134780 84320 1 0 $X=134590 $Y=81360
X798 1 500 497 ICV_7 $T=135700 106080 1 0 $X=135510 $Y=103120
X799 1 506 128 ICV_7 $T=150420 84320 0 0 $X=150230 $Y=84080
X800 1 109 498 ICV_7 $T=152260 78880 0 0 $X=152070 $Y=78640
X801 1 131 508 ICV_7 $T=155940 89760 1 0 $X=155750 $Y=86800
X802 1 130 141 ICV_7 $T=161000 84320 0 0 $X=160810 $Y=84080
X803 1 138 510 ICV_7 $T=161460 122400 1 0 $X=161270 $Y=119440
X804 1 139 503 ICV_7 $T=162380 111520 0 0 $X=162190 $Y=111280
X805 1 144 140 ICV_7 $T=165600 116960 0 0 $X=165410 $Y=116720
X806 1 150 509 ICV_7 $T=175260 116960 0 0 $X=175070 $Y=116720
X807 1 385 3 ICV_7 $T=178020 95200 0 0 $X=177830 $Y=94960
X808 1 109 108 ICV_7 $T=184000 84320 1 0 $X=183810 $Y=81360
X809 1 113 520 ICV_7 $T=184000 89760 1 0 $X=183810 $Y=86800
X810 1 159 4 ICV_7 $T=189520 89760 1 0 $X=189330 $Y=86800
X811 1 522 169 ICV_7 $T=195040 116960 1 0 $X=194850 $Y=114000
X812 1 171 171 ICV_7 $T=197340 122400 1 0 $X=197150 $Y=119440
X813 1 497 8 ICV_7 $T=202400 95200 1 0 $X=202210 $Y=92240
X814 1 528 9 ICV_7 $T=203320 106080 1 0 $X=203130 $Y=103120
X815 1 3 8 ICV_7 $T=203780 100640 1 0 $X=203590 $Y=97680
X816 1 515 530 ICV_7 $T=207000 89760 1 0 $X=206810 $Y=86800
X817 1 160 180 ICV_7 $T=209300 78880 0 0 $X=209110 $Y=78640
X818 1 531 12 ICV_7 $T=212060 95200 0 0 $X=211870 $Y=94960
X819 1 129 183 ICV_7 $T=218040 116960 0 0 $X=217850 $Y=116720
X820 1 133 534 ICV_7 $T=224020 100640 0 0 $X=223830 $Y=100400
X821 1 190 534 ICV_7 $T=224020 106080 0 0 $X=223830 $Y=105840
X822 1 535 189 ICV_7 $T=224480 116960 0 0 $X=224290 $Y=116720
X823 1 536 195 ICV_7 $T=227240 122400 1 0 $X=227050 $Y=119440
X824 1 190 196 ICV_7 $T=228160 116960 1 0 $X=227970 $Y=114000
X825 1 35 40 ICV_7 $T=231380 122400 0 0 $X=231190 $Y=122160
X826 1 208 542 ICV_7 $T=238740 122400 1 0 $X=238550 $Y=119440
X827 1 537 518 ICV_7 $T=240580 89760 0 0 $X=240390 $Y=89520
X828 1 543 211 ICV_7 $T=241960 84320 0 0 $X=241770 $Y=84080
X829 1 12 545 ICV_7 $T=245640 111520 0 0 $X=245450 $Y=111280
X830 1 216 211 ICV_7 $T=250700 84320 0 0 $X=250510 $Y=84080
X831 1 146 219 ICV_7 $T=252540 89760 0 0 $X=252350 $Y=89520
X832 1 549 549 ICV_7 $T=254380 122400 1 0 $X=254190 $Y=119440
X833 1 224 211 ICV_7 $T=258520 84320 1 0 $X=258330 $Y=81360
X834 1 553 225 ICV_7 $T=258520 111520 1 0 $X=258330 $Y=108560
X835 1 555 555 ICV_7 $T=261740 95200 0 0 $X=261550 $Y=94960
X836 1 9 220 ICV_7 $T=264500 89760 0 0 $X=264310 $Y=89520
X837 1 554 229 ICV_7 $T=264500 122400 0 0 $X=264310 $Y=122160
X838 1 226 81 ICV_7 $T=269100 116960 0 0 $X=268910 $Y=116720
X839 1 559 559 ICV_7 $T=273700 95200 1 0 $X=273510 $Y=92240
X840 1 235 221 ICV_7 $T=274620 89760 0 0 $X=274430 $Y=89520
X841 1 564 564 ICV_7 $T=276460 95200 0 0 $X=276270 $Y=94960
X842 1 218 179 ICV_7 $T=280140 116960 0 0 $X=279950 $Y=116720
X843 1 233 220 ICV_7 $T=286120 84320 1 0 $X=285930 $Y=81360
X844 1 566 235 ICV_7 $T=287040 89760 1 0 $X=286850 $Y=86800
X845 1 245 246 ICV_7 $T=292100 95200 0 0 $X=291910 $Y=94960
X846 1 570 198 ICV_7 $T=295320 84320 0 0 $X=295130 $Y=84080
X847 1 572 40 ICV_7 $T=295320 111520 0 0 $X=295130 $Y=111280
X848 1 574 253 ICV_7 $T=298080 106080 0 0 $X=297890 $Y=105840
X849 1 252 49 ICV_7 $T=299000 111520 0 0 $X=298810 $Y=111280
X850 1 527 255 ICV_7 $T=299920 78880 0 0 $X=299730 $Y=78640
X851 1 254 573 ICV_7 $T=300840 122400 0 0 $X=300650 $Y=122160
X852 1 527 240 ICV_7 $T=301300 84320 0 0 $X=301110 $Y=84080
X853 1 167 581 ICV_7 $T=306360 100640 0 0 $X=306170 $Y=100400
X854 1 35 574 ICV_7 $T=308200 106080 0 0 $X=308010 $Y=105840
X855 1 585 12 ICV_7 $T=312340 100640 1 0 $X=312150 $Y=97680
X856 1 167 580 ICV_7 $T=315560 106080 0 0 $X=315370 $Y=105840
X857 1 12 11 ICV_7 $T=324300 89760 0 0 $X=324110 $Y=89520
X858 1 12 11 ICV_7 $T=324300 116960 0 0 $X=324110 $Y=116720
X859 1 11 12 ICV_7 $T=332120 106080 0 0 $X=331930 $Y=105840
X860 1 11 12 ICV_7 $T=333040 95200 0 0 $X=332850 $Y=94960
X861 1 11 12 ICV_7 $T=333040 111520 0 0 $X=332850 $Y=111280
X862 1 11 12 ICV_7 $T=333500 100640 0 0 $X=333310 $Y=100400
X863 1 11 12 ICV_7 $T=334420 78880 0 0 $X=334230 $Y=78640
X864 1 11 12 ICV_7 $T=334880 84320 0 0 $X=334690 $Y=84080
X865 1 2 11 13 12 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 78880 0 0 $X=7630 $Y=78640
X866 1 2 11 14 12 2 19 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 100640 0 0 $X=7630 $Y=100400
X867 1 2 11 15 12 2 20 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 106080 0 0 $X=7630 $Y=105840
X868 1 2 11 16 12 2 21 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 116960 0 0 $X=7630 $Y=116720
X869 1 2 588 406 12 2 23 1 sky130_fd_sc_hd__dfrtp_4 $T=10120 122400 0 0 $X=9930 $Y=122160
X870 1 2 589 407 12 2 26 1 sky130_fd_sc_hd__dfrtp_4 $T=12880 89760 0 0 $X=12690 $Y=89520
X871 1 2 590 409 12 2 27 1 sky130_fd_sc_hd__dfrtp_4 $T=14260 84320 0 0 $X=14070 $Y=84080
X872 1 2 591 417 12 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=23920 122400 1 0 $X=23730 $Y=119440
X873 1 2 592 415 12 2 38 1 sky130_fd_sc_hd__dfrtp_4 $T=27600 84320 1 0 $X=27410 $Y=81360
X874 1 2 593 425 12 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=29900 106080 1 0 $X=29710 $Y=103120
X875 1 2 594 432 12 2 45 1 sky130_fd_sc_hd__dfrtp_4 $T=42320 116960 0 0 $X=42130 $Y=116720
X876 1 2 595 437 12 2 53 1 sky130_fd_sc_hd__dfrtp_4 $T=49220 84320 1 0 $X=49030 $Y=81360
X877 1 2 596 440 12 2 54 1 sky130_fd_sc_hd__dfrtp_4 $T=51060 95200 1 0 $X=50870 $Y=92240
X878 1 2 597 56 12 2 68 1 sky130_fd_sc_hd__dfrtp_4 $T=65780 122400 0 0 $X=65590 $Y=122160
X879 1 2 598 453 12 2 71 1 sky130_fd_sc_hd__dfrtp_4 $T=77280 122400 1 0 $X=77090 $Y=119440
X880 1 2 599 469 12 2 80 1 sky130_fd_sc_hd__dfrtp_4 $T=87860 84320 1 0 $X=87670 $Y=81360
X881 1 2 600 493 12 2 110 1 sky130_fd_sc_hd__dfrtp_4 $T=121440 116960 0 0 $X=121250 $Y=116720
X882 1 2 601 121 12 2 126 1 sky130_fd_sc_hd__dfrtp_4 $T=147200 122400 0 0 $X=147010 $Y=122160
X883 1 2 602 516 12 2 131 1 sky130_fd_sc_hd__dfrtp_4 $T=170200 100640 1 0 $X=170010 $Y=97680
X884 1 2 603 514 12 2 149 1 sky130_fd_sc_hd__dfrtp_4 $T=175260 122400 0 0 $X=175070 $Y=122160
X885 1 2 604 153 12 2 157 1 sky130_fd_sc_hd__dfrtp_4 $T=178020 100640 0 0 $X=177830 $Y=100400
X886 1 2 605 529 12 2 181 1 sky130_fd_sc_hd__dfrtp_4 $T=208380 106080 0 0 $X=208190 $Y=105840
X887 1 2 606 530 12 2 134 1 sky130_fd_sc_hd__dfrtp_4 $T=208840 89760 0 0 $X=208650 $Y=89520
X888 1 2 607 531 12 2 188 1 sky130_fd_sc_hd__dfrtp_4 $T=215740 95200 0 0 $X=215550 $Y=94960
X889 1 2 608 540 12 2 204 1 sky130_fd_sc_hd__dfrtp_4 $T=233220 106080 0 0 $X=233030 $Y=105840
X890 1 2 609 545 12 2 217 1 sky130_fd_sc_hd__dfrtp_4 $T=245640 116960 1 0 $X=245450 $Y=114000
X891 1 2 610 551 12 2 222 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 100640 0 0 $X=259250 $Y=100400
X892 1 2 611 553 12 2 225 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 111520 0 0 $X=259250 $Y=111280
X893 1 2 612 558 12 2 227 1 sky130_fd_sc_hd__dfrtp_4 $T=273700 100640 1 0 $X=273510 $Y=97680
X894 1 2 613 565 12 2 238 1 sky130_fd_sc_hd__dfrtp_4 $T=280140 111520 1 0 $X=279950 $Y=108560
X895 1 2 614 239 12 2 243 1 sky130_fd_sc_hd__dfrtp_4 $T=287500 122400 0 0 $X=287310 $Y=122160
X896 1 2 615 584 12 2 264 1 sky130_fd_sc_hd__dfrtp_4 $T=312340 122400 1 0 $X=312150 $Y=119440
X897 1 2 616 583 12 2 587 1 sky130_fd_sc_hd__dfrtp_4 $T=314180 106080 1 0 $X=313990 $Y=103120
X898 1 2 617 266 12 2 258 1 sky130_fd_sc_hd__dfrtp_4 $T=315560 84320 0 0 $X=315370 $Y=84080
X899 1 2 618 585 12 2 586 1 sky130_fd_sc_hd__dfrtp_4 $T=315560 100640 0 0 $X=315370 $Y=100400
X900 1 2 619 268 12 2 271 1 sky130_fd_sc_hd__dfrtp_4 $T=316940 122400 0 0 $X=316750 $Y=122160
X901 1 2 11 587 12 2 279 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 89760 0 0 $X=327790 $Y=89520
X902 1 2 11 272 12 2 280 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 116960 0 0 $X=327790 $Y=116720
X903 1 2 11 274 12 2 282 1 sky130_fd_sc_hd__dfrtp_4 $T=332120 111520 1 0 $X=331930 $Y=108560
X904 1 2 11 586 12 2 283 1 sky130_fd_sc_hd__dfrtp_4 $T=333040 95200 1 0 $X=332850 $Y=92240
X905 1 2 11 275 12 2 284 1 sky130_fd_sc_hd__dfrtp_4 $T=333040 100640 1 0 $X=332850 $Y=97680
X906 1 2 11 276 12 2 285 1 sky130_fd_sc_hd__dfrtp_4 $T=333040 116960 1 0 $X=332850 $Y=114000
X907 1 2 11 271 12 2 286 1 sky130_fd_sc_hd__dfrtp_4 $T=333500 106080 1 0 $X=333310 $Y=103120
X908 1 2 11 273 12 2 287 1 sky130_fd_sc_hd__dfrtp_4 $T=333960 122400 1 0 $X=333770 $Y=119440
X909 1 2 11 277 12 2 288 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 84320 1 0 $X=334230 $Y=81360
X910 1 2 11 278 12 2 289 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 89760 1 0 $X=334690 $Y=86800
X911 1 2 426 ICV_12 $T=31280 106080 0 0 $X=31090 $Y=105840
X912 1 2 47 ICV_12 $T=50600 100640 1 0 $X=50410 $Y=97680
X913 1 2 444 ICV_12 $T=59800 111520 1 0 $X=59610 $Y=108560
X914 1 2 76 ICV_12 $T=101660 111520 0 0 $X=101470 $Y=111280
X915 1 2 501 ICV_12 $T=147200 95200 0 0 $X=147010 $Y=94960
X916 1 2 143 ICV_12 $T=167900 122400 0 0 $X=167710 $Y=122160
X917 1 2 5 ICV_12 $T=195960 84320 0 0 $X=195770 $Y=84080
X918 1 2 161 ICV_12 $T=199640 95200 0 0 $X=199450 $Y=94960
X919 1 2 532 ICV_12 $T=218960 100640 1 0 $X=218770 $Y=97680
X920 1 2 183 ICV_12 $T=227700 100640 0 0 $X=227510 $Y=100400
X921 1 2 541 ICV_12 $T=241960 116960 1 0 $X=241770 $Y=114000
X922 1 2 550 ICV_12 $T=255760 95200 0 0 $X=255570 $Y=94960
X923 1 2 221 ICV_12 $T=256220 84320 1 0 $X=256030 $Y=81360
X924 1 2 226 ICV_12 $T=266800 116960 0 0 $X=266610 $Y=116720
X925 1 2 222 ICV_12 $T=272320 89760 0 0 $X=272130 $Y=89520
X926 1 2 563 ICV_12 $T=283820 116960 0 0 $X=283630 $Y=116720
X927 1 2 233 ICV_12 $T=284740 89760 1 0 $X=284550 $Y=86800
X928 1 2 569 ICV_12 $T=289800 95200 0 0 $X=289610 $Y=94960
X929 1 2 576 ICV_12 $T=311880 106080 0 0 $X=311690 $Y=105840
X930 1 2 24 ICV_13 $T=19780 95200 0 0 $X=19590 $Y=94960
X931 1 2 25 ICV_13 $T=20240 100640 1 0 $X=20050 $Y=97680
X932 1 2 23 ICV_13 $T=20700 122400 0 0 $X=20510 $Y=122160
X933 1 2 27 ICV_13 $T=23920 84320 1 0 $X=23730 $Y=81360
X934 1 2 31 ICV_13 $T=29900 95200 0 0 $X=29710 $Y=94960
X935 1 2 426 ICV_13 $T=30360 100640 1 0 $X=30170 $Y=97680
X936 1 2 423 ICV_13 $T=32660 116960 1 0 $X=32470 $Y=114000
X937 1 2 36 ICV_13 $T=34500 122400 1 0 $X=34310 $Y=119440
X938 1 2 12 ICV_13 $T=38640 116960 0 0 $X=38450 $Y=116720
X939 1 2 430 ICV_13 $T=43240 106080 0 0 $X=43050 $Y=105840
X940 1 2 438 ICV_13 $T=47380 100640 0 0 $X=47190 $Y=100400
X941 1 2 443 ICV_13 $T=57960 78880 0 0 $X=57770 $Y=78640
X942 1 2 12 ICV_13 $T=62100 122400 0 0 $X=61910 $Y=122160
X943 1 2 59 ICV_13 $T=72220 111520 1 0 $X=72030 $Y=108560
X944 1 2 467 ICV_13 $T=92460 95200 1 0 $X=92270 $Y=92240
X945 1 2 78 ICV_13 $T=94300 116960 0 0 $X=94110 $Y=116720
X946 1 2 472 ICV_13 $T=106260 95200 0 0 $X=106070 $Y=94960
X947 1 2 99 ICV_13 $T=132020 116960 0 0 $X=131830 $Y=116720
X948 1 2 107 ICV_13 $T=141220 100640 1 0 $X=141030 $Y=97680
X949 1 2 501 ICV_13 $T=142600 95200 1 0 $X=142410 $Y=92240
X950 1 2 500 ICV_13 $T=143520 84320 1 0 $X=143330 $Y=81360
X951 1 2 502 ICV_13 $T=143980 89760 1 0 $X=143790 $Y=86800
X952 1 2 498 ICV_13 $T=170200 84320 0 0 $X=170010 $Y=84080
X953 1 2 149 ICV_13 $T=171120 122400 1 0 $X=170930 $Y=119440
X954 1 2 12 ICV_13 $T=174340 100640 0 0 $X=174150 $Y=100400
X955 1 2 518 ICV_13 $T=176180 89760 1 0 $X=175990 $Y=86800
X956 1 2 93 ICV_13 $T=179400 78880 0 0 $X=179210 $Y=78640
X957 1 2 522 ICV_13 $T=190900 111520 0 0 $X=190710 $Y=111280
X958 1 2 519 ICV_13 $T=194580 106080 0 0 $X=194390 $Y=105840
X959 1 2 152 ICV_13 $T=198260 78880 0 0 $X=198070 $Y=78640
X960 1 2 174 ICV_13 $T=198260 116960 0 0 $X=198070 $Y=116720
X961 1 2 173 ICV_13 $T=200100 116960 1 0 $X=199910 $Y=114000
X962 1 2 433 ICV_13 $T=214820 122400 0 0 $X=214630 $Y=122160
X963 1 2 201 ICV_13 $T=233680 78880 0 0 $X=233490 $Y=78640
X964 1 2 197 ICV_13 $T=238280 116960 0 0 $X=238090 $Y=116720
X965 1 2 538 ICV_13 $T=240580 111520 1 0 $X=240390 $Y=108560
X966 1 2 212 ICV_13 $T=242880 78880 0 0 $X=242690 $Y=78640
X967 1 2 544 ICV_13 $T=242880 95200 0 0 $X=242690 $Y=94960
X968 1 2 116 ICV_13 $T=243800 122400 0 0 $X=243610 $Y=122160
X969 1 2 537 ICV_13 $T=244720 100640 1 0 $X=244530 $Y=97680
X970 1 2 214 ICV_13 $T=252540 89760 1 0 $X=252350 $Y=86800
X971 1 2 220 ICV_13 $T=252540 95200 1 0 $X=252350 $Y=92240
X972 1 2 223 ICV_13 $T=254380 116960 0 0 $X=254190 $Y=116720
X973 1 2 169 ICV_13 $T=256220 116960 1 0 $X=256030 $Y=114000
X974 1 2 230 ICV_13 $T=277380 78880 0 0 $X=277190 $Y=78640
X975 1 2 230 ICV_13 $T=282440 78880 0 0 $X=282250 $Y=78640
X976 1 2 221 ICV_13 $T=282440 89760 0 0 $X=282250 $Y=89520
X977 1 2 241 ICV_13 $T=286580 84320 0 0 $X=286390 $Y=84080
X978 1 2 ICV_14 $T=19780 95200 1 0 $X=19590 $Y=92240
X979 1 2 ICV_14 $T=33580 84320 0 0 $X=33390 $Y=84080
X980 1 2 ICV_14 $T=33580 111520 0 0 $X=33390 $Y=111280
X981 1 2 ICV_14 $T=47840 100640 1 0 $X=47650 $Y=97680
X982 1 2 ICV_14 $T=47840 106080 1 0 $X=47650 $Y=103120
X983 1 2 ICV_14 $T=61640 89760 0 0 $X=61450 $Y=89520
X984 1 2 ICV_14 $T=61640 106080 0 0 $X=61450 $Y=105840
X985 1 2 ICV_14 $T=75900 95200 1 0 $X=75710 $Y=92240
X986 1 2 ICV_14 $T=75900 116960 1 0 $X=75710 $Y=114000
X987 1 2 ICV_14 $T=89700 106080 0 0 $X=89510 $Y=105840
X988 1 2 ICV_14 $T=89700 111520 0 0 $X=89510 $Y=111280
X989 1 2 ICV_14 $T=103960 111520 1 0 $X=103770 $Y=108560
X990 1 2 ICV_14 $T=103960 116960 1 0 $X=103770 $Y=114000
X991 1 2 ICV_14 $T=103960 122400 1 0 $X=103770 $Y=119440
X992 1 2 ICV_14 $T=117760 84320 0 0 $X=117570 $Y=84080
X993 1 2 ICV_14 $T=132020 84320 1 0 $X=131830 $Y=81360
X994 1 2 ICV_14 $T=132020 89760 1 0 $X=131830 $Y=86800
X995 1 2 ICV_14 $T=132020 95200 1 0 $X=131830 $Y=92240
X996 1 2 ICV_14 $T=216200 100640 1 0 $X=216010 $Y=97680
X997 1 2 ICV_14 $T=230000 78880 0 0 $X=229810 $Y=78640
X998 1 2 ICV_14 $T=328440 95200 1 0 $X=328250 $Y=92240
X999 1 26 ICV_15 $T=31740 89760 0 0 $X=31550 $Y=89520
X1000 1 426 ICV_15 $T=31740 116960 0 0 $X=31550 $Y=116720
X1001 1 54 ICV_15 $T=59800 95200 0 0 $X=59610 $Y=94960
X1002 1 455 ICV_15 $T=74060 100640 1 0 $X=73870 $Y=97680
X1003 1 12 ICV_15 $T=87860 78880 0 0 $X=87670 $Y=78640
X1004 1 481 ICV_15 $T=102120 100640 1 0 $X=101930 $Y=97680
X1005 1 99 ICV_15 $T=115920 89760 0 0 $X=115730 $Y=89520
X1006 1 100 ICV_15 $T=115920 100640 0 0 $X=115730 $Y=100400
X1007 1 504 ICV_15 $T=143980 89760 0 0 $X=143790 $Y=89520
X1008 1 112 ICV_15 $T=143980 95200 0 0 $X=143790 $Y=94960
X1009 1 12 ICV_15 $T=143980 122400 0 0 $X=143790 $Y=122160
X1010 1 516 ICV_15 $T=172040 95200 0 0 $X=171850 $Y=94960
X1011 1 525 ICV_15 $T=200100 89760 0 0 $X=199910 $Y=89520
X1012 1 184 ICV_15 $T=214360 122400 1 0 $X=214170 $Y=119440
X1013 1 120 ICV_15 $T=228160 116960 0 0 $X=227970 $Y=116720
X1014 1 219 ICV_15 $T=256220 89760 0 0 $X=256030 $Y=89520
X1015 1 12 ICV_15 $T=256220 100640 0 0 $X=256030 $Y=100400
X1016 1 560 ICV_15 $T=270480 116960 1 0 $X=270290 $Y=114000
X1017 1 546 ICV_15 $T=284280 95200 0 0 $X=284090 $Y=94960
X1018 1 238 ICV_15 $T=284280 111520 0 0 $X=284090 $Y=111280
X1019 1 12 ICV_15 $T=284280 122400 0 0 $X=284090 $Y=122160
X1020 1 572 ICV_15 $T=298540 111520 1 0 $X=298350 $Y=108560
X1021 1 575 ICV_15 $T=298540 116960 1 0 $X=298350 $Y=114000
X1022 1 40 ICV_15 $T=298540 122400 1 0 $X=298350 $Y=119440
X1023 1 12 ICV_15 $T=312340 84320 0 0 $X=312150 $Y=84080
X1024 1 2 12 ICV_16 $T=7820 84320 1 0 $X=7630 $Y=81360
X1025 1 2 433 ICV_16 $T=53820 116960 0 0 $X=53630 $Y=116720
X1026 1 2 58 ICV_16 $T=64860 116960 1 0 $X=64670 $Y=114000
X1027 1 2 469 ICV_16 $T=91080 78880 0 0 $X=90890 $Y=78640
X1028 1 2 86 ICV_16 $T=104420 122400 0 0 $X=104230 $Y=122160
X1029 1 2 102 ICV_16 $T=120060 84320 1 0 $X=119870 $Y=81360
X1030 1 2 493 ICV_16 $T=121440 116960 1 0 $X=121250 $Y=114000
X1031 1 2 496 ICV_16 $T=123740 111520 1 0 $X=123550 $Y=108560
X1032 1 2 459 ICV_16 $T=135700 122400 1 0 $X=135510 $Y=119440
X1033 1 2 503 ICV_16 $T=136160 106080 0 0 $X=135970 $Y=105840
X1034 1 2 505 ICV_16 $T=152720 100640 1 0 $X=152530 $Y=97680
X1035 1 2 433 ICV_16 $T=155020 116960 0 0 $X=154830 $Y=116720
X1036 1 2 127 ICV_16 $T=155480 111520 0 0 $X=155290 $Y=111280
X1037 1 2 132 ICV_16 $T=158240 106080 0 0 $X=158050 $Y=105840
X1038 1 2 134 ICV_16 $T=162380 100640 0 0 $X=162190 $Y=100400
X1039 1 2 504 ICV_16 $T=163760 95200 1 0 $X=163570 $Y=92240
X1040 1 2 153 ICV_16 $T=178020 106080 1 0 $X=177830 $Y=103120
X1041 1 2 157 ICV_16 $T=180320 106080 0 0 $X=180130 $Y=105840
X1042 1 2 388 ICV_16 $T=181700 100640 1 0 $X=181510 $Y=97680
X1043 1 2 160 ICV_16 $T=187680 89760 0 0 $X=187490 $Y=89520
X1044 1 2 526 ICV_16 $T=207460 122400 1 0 $X=207270 $Y=119440
X1045 1 2 529 ICV_16 $T=208380 111520 1 0 $X=208190 $Y=108560
X1046 1 2 524 ICV_16 $T=210220 84320 0 0 $X=210030 $Y=84080
X1047 1 2 401 ICV_16 $T=210680 111520 0 0 $X=210490 $Y=111280
X1048 1 2 188 ICV_16 $T=221260 95200 1 0 $X=221070 $Y=92240
X1049 1 2 204 ICV_16 $T=236440 106080 1 0 $X=236250 $Y=103120
X1050 1 2 192 ICV_16 $T=244720 106080 0 0 $X=244530 $Y=105840
X1051 1 2 196 ICV_16 $T=247480 122400 1 0 $X=247290 $Y=119440
X1052 1 2 551 ICV_16 $T=258520 106080 1 0 $X=258330 $Y=103120
X1053 1 2 243 ICV_16 $T=289800 122400 1 0 $X=289610 $Y=119440
X1054 1 2 527 ICV_16 $T=307740 89760 0 0 $X=307550 $Y=89520
X1055 1 2 264 ICV_16 $T=315100 116960 1 0 $X=314910 $Y=114000
X1056 1 2 586 ICV_16 $T=317400 95200 0 0 $X=317210 $Y=94960
X1057 1 2 267 ICV_16 $T=322460 78880 0 0 $X=322270 $Y=78640
X1058 1 2 274 ICV_16 $T=335800 106080 0 0 $X=335610 $Y=105840
X1059 1 2 23 2 423 1 sky130_fd_sc_hd__inv_8 $T=24380 122400 0 0 $X=24190 $Y=122160
X1060 1 2 27 2 419 1 sky130_fd_sc_hd__inv_8 $T=25760 78880 0 0 $X=25570 $Y=78640
X1061 1 2 29 2 418 1 sky130_fd_sc_hd__inv_8 $T=30360 89760 1 0 $X=30170 $Y=86800
X1062 1 2 26 2 413 1 sky130_fd_sc_hd__inv_8 $T=34960 89760 0 0 $X=34770 $Y=89520
X1063 1 2 32 2 422 1 sky130_fd_sc_hd__inv_8 $T=34960 122400 0 0 $X=34770 $Y=122160
X1064 1 2 38 2 429 1 sky130_fd_sc_hd__inv_8 $T=38640 89760 1 0 $X=38450 $Y=86800
X1065 1 2 37 2 430 1 sky130_fd_sc_hd__inv_8 $T=39100 106080 0 0 $X=38910 $Y=105840
X1066 1 2 45 2 51 1 sky130_fd_sc_hd__inv_8 $T=51060 122400 0 0 $X=50870 $Y=122160
X1067 1 2 53 2 61 1 sky130_fd_sc_hd__inv_8 $T=63020 84320 0 0 $X=62830 $Y=84080
X1068 1 2 54 2 44 1 sky130_fd_sc_hd__inv_8 $T=63020 95200 0 0 $X=62830 $Y=94960
X1069 1 2 71 2 66 1 sky130_fd_sc_hd__inv_8 $T=81420 122400 0 0 $X=81230 $Y=122160
X1070 1 2 80 2 479 1 sky130_fd_sc_hd__inv_8 $T=97060 84320 0 0 $X=96870 $Y=84080
X1071 1 2 110 2 491 1 sky130_fd_sc_hd__inv_8 $T=133400 116960 1 0 $X=133210 $Y=114000
X1072 1 2 134 2 115 1 sky130_fd_sc_hd__inv_8 $T=157320 100640 0 0 $X=157130 $Y=100400
X1073 1 2 128 2 506 1 sky130_fd_sc_hd__inv_8 $T=161460 84320 1 0 $X=161270 $Y=81360
X1074 1 2 130 2 508 1 sky130_fd_sc_hd__inv_8 $T=161460 89760 1 0 $X=161270 $Y=86800
X1075 1 2 131 2 507 1 sky130_fd_sc_hd__inv_8 $T=161460 100640 1 0 $X=161270 $Y=97680
X1076 1 2 157 2 139 1 sky130_fd_sc_hd__inv_8 $T=180320 111520 1 0 $X=180130 $Y=108560
X1077 1 2 156 2 522 1 sky130_fd_sc_hd__inv_8 $T=191820 95200 0 0 $X=191630 $Y=94960
X1078 1 2 145 2 159 1 sky130_fd_sc_hd__inv_8 $T=203320 78880 0 0 $X=203130 $Y=78640
X1079 1 2 181 2 392 1 sky130_fd_sc_hd__inv_8 $T=208380 106080 1 0 $X=208190 $Y=103120
X1080 1 2 188 2 534 1 sky130_fd_sc_hd__inv_8 $T=221260 100640 1 0 $X=221070 $Y=97680
X1081 1 2 537 2 4 1 sky130_fd_sc_hd__inv_8 $T=231380 84320 0 0 $X=231190 $Y=84080
X1082 1 2 201 2 202 1 sky130_fd_sc_hd__inv_8 $T=236440 84320 1 0 $X=236250 $Y=81360
X1083 1 2 204 2 536 1 sky130_fd_sc_hd__inv_8 $T=236440 111520 1 0 $X=236250 $Y=108560
X1084 1 2 543 2 191 1 sky130_fd_sc_hd__inv_8 $T=246100 89760 0 0 $X=245910 $Y=89520
X1085 1 2 212 2 214 1 sky130_fd_sc_hd__inv_8 $T=246560 78880 0 0 $X=246370 $Y=78640
X1086 1 2 217 2 208 1 sky130_fd_sc_hd__inv_8 $T=250240 116960 0 0 $X=250050 $Y=116720
X1087 1 2 225 2 549 1 sky130_fd_sc_hd__inv_8 $T=259900 116960 1 0 $X=259710 $Y=114000
X1088 1 2 555 2 547 1 sky130_fd_sc_hd__inv_8 $T=261740 100640 1 0 $X=261550 $Y=97680
X1089 1 2 227 2 548 1 sky130_fd_sc_hd__inv_8 $T=266340 84320 0 0 $X=266150 $Y=84080
X1090 1 2 233 2 564 1 sky130_fd_sc_hd__inv_8 $T=279220 95200 1 0 $X=279030 $Y=92240
X1091 1 2 238 2 560 1 sky130_fd_sc_hd__inv_8 $T=287500 111520 0 0 $X=287310 $Y=111280
X1092 1 2 258 2 262 1 sky130_fd_sc_hd__inv_8 $T=311880 89760 1 0 $X=311690 $Y=86800
X1093 1 2 264 2 573 1 sky130_fd_sc_hd__inv_8 $T=315560 116960 0 0 $X=315370 $Y=116720
X1094 1 2 586 2 572 1 sky130_fd_sc_hd__inv_8 $T=317400 100640 1 0 $X=317210 $Y=97680
X1095 1 2 587 2 574 1 sky130_fd_sc_hd__inv_8 $T=319700 106080 0 0 $X=319510 $Y=105840
X1096 1 2 17 408 2 407 1 sky130_fd_sc_hd__nor2_4 $T=11960 95200 1 0 $X=11770 $Y=92240
X1097 1 2 17 410 2 22 1 sky130_fd_sc_hd__nor2_4 $T=15640 95200 0 0 $X=15450 $Y=94960
X1098 1 2 17 414 2 409 1 sky130_fd_sc_hd__nor2_4 $T=21160 89760 1 0 $X=20970 $Y=86800
X1099 1 2 17 411 2 417 1 sky130_fd_sc_hd__nor2_4 $T=21160 111520 0 0 $X=20970 $Y=111280
X1100 1 2 17 412 2 406 1 sky130_fd_sc_hd__nor2_4 $T=21160 116960 0 0 $X=20970 $Y=116720
X1101 1 2 41 427 2 415 1 sky130_fd_sc_hd__nor2_4 $T=39560 84320 0 0 $X=39370 $Y=84080
X1102 1 2 41 431 2 425 1 sky130_fd_sc_hd__nor2_4 $T=43240 100640 0 0 $X=43050 $Y=100400
X1103 1 2 41 442 2 440 1 sky130_fd_sc_hd__nor2_4 $T=48760 84320 0 0 $X=48570 $Y=84080
X1104 1 2 41 441 2 432 1 sky130_fd_sc_hd__nor2_4 $T=49220 111520 0 0 $X=49030 $Y=111280
X1105 1 2 41 444 2 56 1 sky130_fd_sc_hd__nor2_4 $T=59800 116960 1 0 $X=59610 $Y=114000
X1106 1 2 57 55 2 437 1 sky130_fd_sc_hd__nor2_4 $T=63020 78880 0 0 $X=62830 $Y=78640
X1107 1 2 57 452 2 453 1 sky130_fd_sc_hd__nor2_4 $T=68080 106080 1 0 $X=67890 $Y=103120
X1108 1 2 69 458 2 443 1 sky130_fd_sc_hd__nor2_4 $T=77280 84320 1 0 $X=77090 $Y=81360
X1109 1 2 460 463 2 451 1 sky130_fd_sc_hd__nor2_4 $T=78660 95200 1 0 $X=78470 $Y=92240
X1110 1 2 460 464 2 449 1 sky130_fd_sc_hd__nor2_4 $T=78660 100640 1 0 $X=78470 $Y=97680
X1111 1 2 460 466 2 457 1 sky130_fd_sc_hd__nor2_4 $T=81880 106080 1 0 $X=81690 $Y=103120
X1112 1 2 460 467 2 456 1 sky130_fd_sc_hd__nor2_4 $T=86480 100640 1 0 $X=86290 $Y=97680
X1113 1 2 460 472 2 455 1 sky130_fd_sc_hd__nor2_4 $T=91080 95200 0 0 $X=90890 $Y=94960
X1114 1 2 77 473 2 79 1 sky130_fd_sc_hd__nor2_4 $T=93380 122400 1 0 $X=93190 $Y=119440
X1115 1 2 77 471 2 469 1 sky130_fd_sc_hd__nor2_4 $T=93840 89760 1 0 $X=93650 $Y=86800
X1116 1 2 77 470 2 82 1 sky130_fd_sc_hd__nor2_4 $T=94760 122400 0 0 $X=94570 $Y=122160
X1117 1 2 458 83 2 477 1 sky130_fd_sc_hd__nor2_4 $T=96140 95200 1 0 $X=95950 $Y=92240
X1118 1 2 464 83 2 482 1 sky130_fd_sc_hd__nor2_4 $T=102580 100640 0 0 $X=102390 $Y=100400
X1119 1 2 463 83 2 481 1 sky130_fd_sc_hd__nor2_4 $T=103500 89760 0 0 $X=103310 $Y=89520
X1120 1 2 85 89 2 88 1 sky130_fd_sc_hd__nor2_4 $T=105340 78880 0 0 $X=105150 $Y=78640
X1121 1 2 77 486 2 92 1 sky130_fd_sc_hd__nor2_4 $T=106720 122400 1 0 $X=106530 $Y=119440
X1122 1 2 466 83 2 487 1 sky130_fd_sc_hd__nor2_4 $T=108560 106080 1 0 $X=108370 $Y=103120
X1123 1 2 96 485 2 91 1 sky130_fd_sc_hd__nor2_4 $T=109940 116960 0 0 $X=109750 $Y=116720
X1124 1 2 467 100 2 490 1 sky130_fd_sc_hd__nor2_4 $T=118680 106080 1 0 $X=118490 $Y=103120
X1125 1 2 96 496 2 493 1 sky130_fd_sc_hd__nor2_4 $T=121900 106080 0 0 $X=121710 $Y=105840
X1126 1 2 472 100 2 489 1 sky130_fd_sc_hd__nor2_4 $T=122820 100640 1 0 $X=122630 $Y=97680
X1127 1 2 89 100 2 492 1 sky130_fd_sc_hd__nor2_4 $T=123280 89760 1 0 $X=123090 $Y=86800
X1128 1 2 150 509 2 514 1 sky130_fd_sc_hd__nor2_4 $T=174800 122400 1 0 $X=174610 $Y=119440
X1129 1 2 167 528 2 529 1 sky130_fd_sc_hd__nor2_4 $T=203320 111520 1 0 $X=203130 $Y=108560
X1130 1 2 179 178 2 163 1 sky130_fd_sc_hd__nor2_4 $T=203320 122400 0 0 $X=203130 $Y=122160
X1131 1 2 185 532 2 531 1 sky130_fd_sc_hd__nor2_4 $T=218960 100640 0 0 $X=218770 $Y=100400
X1132 1 2 521 537 2 165 1 sky130_fd_sc_hd__nor2_4 $T=231840 100640 1 0 $X=231650 $Y=97680
X1133 1 2 197 539 2 540 1 sky130_fd_sc_hd__nor2_4 $T=231840 116960 1 0 $X=231650 $Y=114000
X1134 1 2 537 206 2 203 1 sky130_fd_sc_hd__nor2_4 $T=236440 95200 1 0 $X=236250 $Y=92240
X1135 1 2 537 207 2 210 1 sky130_fd_sc_hd__nor2_4 $T=238740 95200 0 0 $X=238550 $Y=94960
X1136 1 2 197 541 2 545 1 sky130_fd_sc_hd__nor2_4 $T=241960 116960 0 0 $X=241770 $Y=116720
X1137 1 2 537 544 2 538 1 sky130_fd_sc_hd__nor2_4 $T=246560 95200 0 0 $X=246370 $Y=94960
X1138 1 2 179 554 2 553 1 sky130_fd_sc_hd__nor2_4 $T=259440 122400 0 0 $X=259250 $Y=122160
X1139 1 2 179 562 2 565 1 sky130_fd_sc_hd__nor2_4 $T=275540 116960 1 0 $X=275350 $Y=114000
X1140 1 2 179 563 2 239 1 sky130_fd_sc_hd__nor2_4 $T=281980 122400 1 0 $X=281790 $Y=119440
X1141 1 2 198 237 2 246 1 sky130_fd_sc_hd__nor2_4 $T=290260 84320 1 0 $X=290070 $Y=81360
X1142 1 2 198 241 2 245 1 sky130_fd_sc_hd__nor2_4 $T=290260 84320 0 0 $X=290070 $Y=84080
X1143 1 2 198 570 2 571 1 sky130_fd_sc_hd__nor2_4 $T=291180 89760 1 0 $X=290990 $Y=86800
X1144 1 2 546 245 2 247 1 sky130_fd_sc_hd__nor2_4 $T=292560 100640 1 0 $X=292370 $Y=97680
X1145 1 2 546 571 2 249 1 sky130_fd_sc_hd__nor2_4 $T=294860 100640 0 0 $X=294670 $Y=100400
X1146 1 2 546 246 2 250 1 sky130_fd_sc_hd__nor2_4 $T=295780 95200 0 0 $X=295590 $Y=94960
X1147 1 2 167 581 2 583 1 sky130_fd_sc_hd__nor2_4 $T=306360 106080 1 0 $X=306170 $Y=103120
X1148 1 2 167 578 2 584 1 sky130_fd_sc_hd__nor2_4 $T=310040 116960 1 0 $X=309850 $Y=114000
X1149 1 2 167 580 2 585 1 sky130_fd_sc_hd__nor2_4 $T=314180 111520 1 0 $X=313990 $Y=108560
X1150 1 2 418 25 24 421 2 410 1 sky130_fd_sc_hd__o22a_4 $T=23460 95200 0 0 $X=23270 $Y=94960
X1151 1 2 413 25 24 416 2 408 1 sky130_fd_sc_hd__o22a_4 $T=23920 100640 1 0 $X=23730 $Y=97680
X1152 1 2 419 25 24 424 2 414 1 sky130_fd_sc_hd__o22a_4 $T=24380 95200 1 0 $X=24190 $Y=92240
X1153 1 2 422 25 24 420 2 411 1 sky130_fd_sc_hd__o22a_4 $T=26220 116960 1 0 $X=26030 $Y=114000
X1154 1 2 423 40 35 428 2 412 1 sky130_fd_sc_hd__o22a_4 $T=36340 116960 1 0 $X=36150 $Y=114000
X1155 1 2 44 46 52 434 2 442 1 sky130_fd_sc_hd__o22a_4 $T=51520 78880 0 0 $X=51330 $Y=78640
X1156 1 2 429 46 439 436 2 427 1 sky130_fd_sc_hd__o22a_4 $T=51520 89760 0 0 $X=51330 $Y=89520
X1157 1 2 430 46 439 435 2 431 1 sky130_fd_sc_hd__o22a_4 $T=52900 100640 1 0 $X=52710 $Y=97680
X1158 1 2 51 58 439 448 2 441 1 sky130_fd_sc_hd__o22a_4 $T=63020 111520 0 0 $X=62830 $Y=111280
X1159 1 2 60 64 44 443 2 434 1 sky130_fd_sc_hd__o22a_4 $T=64400 84320 1 0 $X=64210 $Y=81360
X1160 1 2 445 446 429 451 2 436 1 sky130_fd_sc_hd__o22a_4 $T=65780 95200 1 0 $X=65590 $Y=92240
X1161 1 2 59 58 439 447 2 444 1 sky130_fd_sc_hd__o22a_4 $T=65780 111520 1 0 $X=65590 $Y=108560
X1162 1 2 445 450 430 449 2 435 1 sky130_fd_sc_hd__o22a_4 $T=66700 100640 0 0 $X=66510 $Y=100400
X1163 1 2 66 58 439 454 2 452 1 sky130_fd_sc_hd__o22a_4 $T=69460 106080 0 0 $X=69270 $Y=105840
X1164 1 2 445 462 59 456 2 447 1 sky130_fd_sc_hd__o22a_4 $T=77280 111520 1 0 $X=77090 $Y=108560
X1165 1 2 445 465 66 455 2 454 1 sky130_fd_sc_hd__o22a_4 $T=78660 100640 0 0 $X=78470 $Y=100400
X1166 1 2 445 461 51 457 2 448 1 sky130_fd_sc_hd__o22a_4 $T=79580 106080 0 0 $X=79390 $Y=105840
X1167 1 2 64 476 76 477 2 474 1 sky130_fd_sc_hd__o22a_4 $T=93840 106080 1 0 $X=93650 $Y=103120
X1168 1 2 76 78 475 474 2 473 1 sky130_fd_sc_hd__o22a_4 $T=94300 111520 0 0 $X=94110 $Y=111280
X1169 1 2 84 78 475 478 2 470 1 sky130_fd_sc_hd__o22a_4 $T=97980 116960 0 0 $X=97790 $Y=116720
X1170 1 2 450 476 84 482 2 478 1 sky130_fd_sc_hd__o22a_4 $T=98900 106080 0 0 $X=98710 $Y=105840
X1171 1 2 446 476 479 481 2 480 1 sky130_fd_sc_hd__o22a_4 $T=99820 95200 0 0 $X=99630 $Y=94960
X1172 1 2 479 483 475 480 2 471 1 sky130_fd_sc_hd__o22a_4 $T=105340 95200 1 0 $X=105150 $Y=92240
X1173 1 2 461 476 94 487 2 484 1 sky130_fd_sc_hd__o22a_4 $T=106260 111520 1 0 $X=106070 $Y=108560
X1174 1 2 95 483 475 488 2 485 1 sky130_fd_sc_hd__o22a_4 $T=107640 111520 0 0 $X=107450 $Y=111280
X1175 1 2 94 483 475 484 2 486 1 sky130_fd_sc_hd__o22a_4 $T=108560 116960 1 0 $X=108370 $Y=114000
X1176 1 2 462 476 95 490 2 488 1 sky130_fd_sc_hd__o22a_4 $T=116380 111520 1 0 $X=116190 $Y=108560
X1177 1 2 465 101 99 489 2 494 1 sky130_fd_sc_hd__o22a_4 $T=120980 95200 1 0 $X=120790 $Y=92240
X1178 1 2 97 101 491 492 2 495 1 sky130_fd_sc_hd__o22a_4 $T=120980 95200 0 0 $X=120790 $Y=94960
X1179 1 2 99 483 103 494 2 104 1 sky130_fd_sc_hd__o22a_4 $T=122820 89760 0 0 $X=122630 $Y=89520
X1180 1 2 491 483 103 495 2 496 1 sky130_fd_sc_hd__o22a_4 $T=122820 100640 0 0 $X=122630 $Y=100400
X1181 1 2 140 138 135 510 2 509 1 sky130_fd_sc_hd__o22a_4 $T=160540 122400 0 0 $X=160350 $Y=122160
X1182 1 2 392 166 175 401 2 528 1 sky130_fd_sc_hd__o22a_4 $T=203320 111520 0 0 $X=203130 $Y=111280
X1183 1 2 171 173 177 526 2 178 1 sky130_fd_sc_hd__o22a_4 $T=203320 116960 0 0 $X=203130 $Y=116720
X1184 1 2 184 36 433 186 2 187 1 sky130_fd_sc_hd__o22a_4 $T=218500 122400 0 0 $X=218310 $Y=122160
X1185 1 2 534 190 189 533 2 532 1 sky130_fd_sc_hd__o22a_4 $T=222180 111520 1 0 $X=221990 $Y=108560
X1186 1 2 536 190 189 535 2 539 1 sky130_fd_sc_hd__o22a_4 $T=231840 116960 0 0 $X=231650 $Y=116720
X1187 1 2 208 190 189 542 2 541 1 sky130_fd_sc_hd__o22a_4 $T=237360 122400 0 0 $X=237170 $Y=122160
X1188 1 2 549 218 226 552 2 554 1 sky130_fd_sc_hd__o22a_4 $T=259440 116960 0 0 $X=259250 $Y=116720
X1189 1 2 560 218 226 561 2 562 1 sky130_fd_sc_hd__o22a_4 $T=272780 116960 0 0 $X=272590 $Y=116720
X1190 1 2 231 218 226 236 2 563 1 sky130_fd_sc_hd__o22a_4 $T=274160 122400 0 0 $X=273970 $Y=122160
X1191 1 2 573 40 35 575 2 578 1 sky130_fd_sc_hd__o22a_4 $T=302680 116960 0 0 $X=302490 $Y=116720
X1192 1 2 572 40 35 577 2 580 1 sky130_fd_sc_hd__o22a_4 $T=303140 111520 0 0 $X=302950 $Y=111280
X1193 1 2 574 40 35 576 2 581 1 sky130_fd_sc_hd__o22a_4 $T=304060 111520 1 0 $X=303870 $Y=108560
X1194 1 2 36 2 25 1 sky130_fd_sc_hd__buf_1 $T=37260 116960 0 0 $X=37070 $Y=116720
X1195 1 2 433 2 24 1 sky130_fd_sc_hd__buf_1 $T=44160 111520 0 0 $X=43970 $Y=111280
X1196 1 2 42 2 426 1 sky130_fd_sc_hd__buf_1 $T=45540 122400 0 0 $X=45350 $Y=122160
X1197 1 2 36 2 40 1 sky130_fd_sc_hd__buf_1 $T=51060 116960 1 0 $X=50870 $Y=114000
X1198 1 2 433 2 35 1 sky130_fd_sc_hd__buf_1 $T=51980 122400 1 0 $X=51790 $Y=119440
X1199 1 2 70 2 445 1 sky130_fd_sc_hd__buf_1 $T=77740 84320 0 0 $X=77550 $Y=84080
X1200 1 2 459 2 50 1 sky130_fd_sc_hd__buf_1 $T=78660 116960 1 0 $X=78470 $Y=114000
X1201 1 2 72 2 460 1 sky130_fd_sc_hd__buf_1 $T=84180 78880 0 0 $X=83990 $Y=78640
X1202 1 2 459 2 75 1 sky130_fd_sc_hd__buf_1 $T=88320 111520 1 0 $X=88130 $Y=108560
X1203 1 2 459 2 73 1 sky130_fd_sc_hd__buf_1 $T=97060 89760 0 0 $X=96870 $Y=89520
X1204 1 2 93 2 483 1 sky130_fd_sc_hd__buf_1 $T=110860 89760 1 0 $X=110670 $Y=86800
X1205 1 2 98 2 475 1 sky130_fd_sc_hd__buf_1 $T=115920 89760 1 0 $X=115730 $Y=86800
X1206 1 2 102 2 476 1 sky130_fd_sc_hd__buf_1 $T=120060 84320 0 0 $X=119870 $Y=84080
X1207 1 2 459 2 105 1 sky130_fd_sc_hd__buf_1 $T=133400 122400 1 0 $X=133210 $Y=119440
X1208 1 2 503 2 438 1 sky130_fd_sc_hd__buf_1 $T=136160 111520 1 0 $X=135970 $Y=108560
X1209 1 2 112 2 111 1 sky130_fd_sc_hd__buf_1 $T=144900 100640 1 0 $X=144710 $Y=97680
X1210 1 2 502 2 498 1 sky130_fd_sc_hd__buf_1 $T=147200 84320 0 0 $X=147010 $Y=84080
X1211 1 2 500 2 109 1 sky130_fd_sc_hd__buf_1 $T=147660 89760 1 0 $X=147470 $Y=86800
X1212 1 2 115 2 497 1 sky130_fd_sc_hd__buf_1 $T=149500 95200 0 0 $X=149310 $Y=94960
X1213 1 2 505 2 464 1 sky130_fd_sc_hd__buf_1 $T=150420 100640 1 0 $X=150230 $Y=97680
X1214 1 2 506 2 107 1 sky130_fd_sc_hd__buf_1 $T=152720 89760 1 0 $X=152530 $Y=86800
X1215 1 2 508 2 501 1 sky130_fd_sc_hd__buf_1 $T=154100 95200 1 0 $X=153910 $Y=92240
X1216 1 2 131 2 502 1 sky130_fd_sc_hd__buf_1 $T=154560 95200 0 0 $X=154370 $Y=94960
X1217 1 2 107 2 108 1 sky130_fd_sc_hd__buf_1 $T=155020 84320 1 0 $X=154830 $Y=81360
X1218 1 2 433 2 135 1 sky130_fd_sc_hd__buf_1 $T=155020 122400 1 0 $X=154830 $Y=119440
X1219 1 2 504 2 114 1 sky130_fd_sc_hd__buf_1 $T=161460 95200 1 0 $X=161270 $Y=92240
X1220 1 2 134 2 504 1 sky130_fd_sc_hd__buf_1 $T=161460 106080 1 0 $X=161270 $Y=103120
X1221 1 2 130 2 499 1 sky130_fd_sc_hd__buf_1 $T=163300 89760 0 0 $X=163110 $Y=89520
X1222 1 2 511 2 503 1 sky130_fd_sc_hd__buf_1 $T=164680 111520 1 0 $X=164490 $Y=108560
X1223 1 2 158 2 150 1 sky130_fd_sc_hd__buf_1 $T=183080 122400 1 0 $X=182890 $Y=119440
X1224 1 2 161 2 519 1 sky130_fd_sc_hd__buf_1 $T=189520 111520 1 0 $X=189330 $Y=108560
X1225 1 2 42 2 147 1 sky130_fd_sc_hd__buf_1 $T=189520 122400 1 0 $X=189330 $Y=119440
X1226 1 2 165 2 166 1 sky130_fd_sc_hd__buf_1 $T=193660 122400 1 0 $X=193470 $Y=119440
X1227 1 2 156 2 9 1 sky130_fd_sc_hd__buf_1 $T=194580 95200 1 0 $X=194390 $Y=92240
X1228 1 2 522 2 161 1 sky130_fd_sc_hd__buf_1 $T=194580 111520 0 0 $X=194390 $Y=111280
X1229 1 2 519 2 168 1 sky130_fd_sc_hd__buf_1 $T=196420 111520 1 0 $X=196230 $Y=108560
X1230 1 2 522 2 170 1 sky130_fd_sc_hd__buf_1 $T=196880 116960 0 0 $X=196690 $Y=116720
X1231 1 2 36 2 173 1 sky130_fd_sc_hd__buf_1 $T=198720 116960 1 0 $X=198530 $Y=114000
X1232 1 2 525 2 145 1 sky130_fd_sc_hd__buf_1 $T=203320 89760 0 0 $X=203130 $Y=89520
X1233 1 2 182 2 183 1 sky130_fd_sc_hd__buf_1 $T=213440 122400 0 0 $X=213250 $Y=122160
X1234 1 2 158 2 185 1 sky130_fd_sc_hd__buf_1 $T=214820 116960 0 0 $X=214630 $Y=116720
X1235 1 2 191 2 433 1 sky130_fd_sc_hd__buf_1 $T=224940 111520 0 0 $X=224750 $Y=111280
X1236 1 2 192 2 194 1 sky130_fd_sc_hd__buf_1 $T=228620 84320 1 0 $X=228430 $Y=81360
X1237 1 2 198 2 152 1 sky130_fd_sc_hd__buf_1 $T=232300 78880 0 0 $X=232110 $Y=78640
X1238 1 2 199 2 200 1 sky130_fd_sc_hd__buf_1 $T=234140 89760 1 0 $X=233950 $Y=86800
X1239 1 2 191 2 189 1 sky130_fd_sc_hd__buf_1 $T=237360 111520 0 0 $X=237170 $Y=111280
X1240 1 2 538 2 190 1 sky130_fd_sc_hd__buf_1 $T=242420 111520 0 0 $X=242230 $Y=111280
X1241 1 2 518 2 546 1 sky130_fd_sc_hd__buf_1 $T=245640 95200 1 0 $X=245450 $Y=92240
X1242 1 2 192 2 215 1 sky130_fd_sc_hd__buf_1 $T=245640 111520 1 0 $X=245450 $Y=108560
X1243 1 2 538 2 218 1 sky130_fd_sc_hd__buf_1 $T=251620 111520 0 0 $X=251430 $Y=111280
X1244 1 2 557 2 212 1 sky130_fd_sc_hd__buf_1 $T=263120 89760 1 0 $X=262930 $Y=86800
X1245 1 2 556 2 555 1 sky130_fd_sc_hd__buf_1 $T=265420 95200 1 0 $X=265230 $Y=92240
X1246 1 2 222 2 233 1 sky130_fd_sc_hd__buf_1 $T=270020 89760 0 0 $X=269830 $Y=89520
X1247 1 2 221 2 219 1 sky130_fd_sc_hd__buf_1 $T=273700 84320 1 0 $X=273510 $Y=81360
X1248 1 2 191 2 226 1 sky130_fd_sc_hd__buf_1 $T=276920 111520 0 0 $X=276730 $Y=111280
X1249 1 2 564 2 220 1 sky130_fd_sc_hd__buf_1 $T=280600 95200 0 0 $X=280410 $Y=94960
X1250 1 2 235 2 198 1 sky130_fd_sc_hd__buf_1 $T=281060 78880 0 0 $X=280870 $Y=78640
X1251 1 2 566 2 240 1 sky130_fd_sc_hd__buf_1 $T=287040 95200 1 0 $X=286850 $Y=92240
X1252 1 2 546 2 8 1 sky130_fd_sc_hd__buf_1 $T=287040 100640 1 0 $X=286850 $Y=97680
X1253 1 2 569 2 242 1 sky130_fd_sc_hd__buf_1 $T=287500 95200 0 0 $X=287310 $Y=94960
X1254 1 2 28 422 426 2 420 1 sky130_fd_sc_hd__o21a_4 $T=29440 111520 1 0 $X=29250 $Y=108560
X1255 1 2 33 418 426 2 421 1 sky130_fd_sc_hd__o21a_4 $T=34040 100640 1 0 $X=33850 $Y=97680
X1256 1 2 31 419 426 2 424 1 sky130_fd_sc_hd__o21a_4 $T=34960 95200 0 0 $X=34770 $Y=94960
X1257 1 2 39 413 426 2 416 1 sky130_fd_sc_hd__o21a_4 $T=34960 100640 0 0 $X=34770 $Y=100400
X1258 1 2 34 423 426 2 428 1 sky130_fd_sc_hd__o21a_4 $T=38180 122400 1 0 $X=37990 $Y=119440
X1259 1 2 141 464 145 2 142 1 sky130_fd_sc_hd__o21a_4 $T=164680 84320 0 0 $X=164490 $Y=84080
X1260 1 2 144 140 147 2 510 1 sky130_fd_sc_hd__o21a_4 $T=165600 122400 1 0 $X=165410 $Y=119440
X1261 1 2 148 517 513 2 516 1 sky130_fd_sc_hd__o21a_4 $T=175260 89760 0 0 $X=175070 $Y=89520
X1262 1 2 521 157 519 2 385 1 sky130_fd_sc_hd__o21a_4 $T=189980 100640 1 0 $X=189790 $Y=97680
X1263 1 2 174 171 169 2 526 1 sky130_fd_sc_hd__o21a_4 $T=201020 122400 1 0 $X=200830 $Y=119440
X1264 1 2 129 184 183 2 186 1 sky130_fd_sc_hd__o21a_4 $T=218040 122400 1 0 $X=217850 $Y=119440
X1265 1 2 133 534 183 2 533 1 sky130_fd_sc_hd__o21a_4 $T=223100 106080 1 0 $X=222910 $Y=103120
X1266 1 2 120 536 196 2 535 1 sky130_fd_sc_hd__o21a_4 $T=232300 122400 1 0 $X=232110 $Y=119440
X1267 1 2 4 198 209 2 205 1 sky130_fd_sc_hd__o21a_4 $T=237360 78880 0 0 $X=237170 $Y=78640
X1268 1 2 116 208 196 2 542 1 sky130_fd_sc_hd__o21a_4 $T=247480 122400 0 0 $X=247290 $Y=122160
X1269 1 2 220 219 146 2 550 1 sky130_fd_sc_hd__o21a_4 $T=256220 95200 1 0 $X=256030 $Y=92240
X1270 1 2 223 549 169 2 552 1 sky130_fd_sc_hd__o21a_4 $T=258060 122400 1 0 $X=257870 $Y=119440
X1271 1 2 81 560 169 2 561 1 sky130_fd_sc_hd__o21a_4 $T=273700 122400 1 0 $X=273510 $Y=119440
X1272 1 2 253 574 252 2 576 1 sky130_fd_sc_hd__o21a_4 $T=301760 106080 0 0 $X=301570 $Y=105840
X1273 1 2 49 572 252 2 577 1 sky130_fd_sc_hd__o21a_4 $T=301760 116960 1 0 $X=301570 $Y=114000
X1274 1 2 254 573 252 2 575 1 sky130_fd_sc_hd__o21a_4 $T=301760 122400 1 0 $X=301570 $Y=119440
X1275 1 2 418 33 ICV_21 $T=30820 95200 1 0 $X=30630 $Y=92240
X1276 1 2 434 437 ICV_21 $T=43240 78880 0 0 $X=43050 $Y=78640
X1277 1 2 43 438 ICV_21 $T=43700 84320 0 0 $X=43510 $Y=84080
X1278 1 2 436 440 ICV_21 $T=44620 89760 0 0 $X=44430 $Y=89520
X1279 1 2 69 458 ICV_21 $T=74980 78880 0 0 $X=74790 $Y=78640
X1280 1 2 457 445 ICV_21 $T=76360 106080 1 0 $X=76170 $Y=103120
X1281 1 2 468 468 ICV_21 $T=87860 89760 1 0 $X=87670 $Y=86800
X1282 1 2 471 77 ICV_21 $T=90160 84320 0 0 $X=89970 $Y=84080
X1283 1 2 473 77 ICV_21 $T=90160 116960 0 0 $X=89970 $Y=116720
X1284 1 2 107 498 ICV_21 $T=127420 78880 0 0 $X=127230 $Y=78640
X1285 1 2 497 497 ICV_21 $T=127420 95200 0 0 $X=127230 $Y=94960
X1286 1 2 107 500 ICV_21 $T=129260 89760 0 0 $X=129070 $Y=89520
X1287 1 2 151 152 ICV_21 $T=174340 84320 0 0 $X=174150 $Y=84080
X1288 1 2 113 5 ICV_21 $T=187220 78880 0 0 $X=187030 $Y=78640
X1289 1 2 519 156 ICV_21 $T=188600 95200 1 0 $X=188410 $Y=92240
X1290 1 2 533 189 ICV_21 $T=218960 106080 0 0 $X=218770 $Y=105840
X1291 1 2 521 537 ICV_21 $T=230460 95200 0 0 $X=230270 $Y=94960
X1292 1 2 215 547 ICV_21 $T=250700 95200 0 0 $X=250510 $Y=94960
X1293 1 2 179 179 ICV_21 $T=253000 122400 0 0 $X=252810 $Y=122160
X1294 1 2 231 169 ICV_21 $T=267260 122400 0 0 $X=267070 $Y=122160
X1295 1 2 12 558 ICV_21 $T=271400 95200 0 0 $X=271210 $Y=94960
X1296 1 2 12 565 ICV_21 $T=278760 106080 0 0 $X=278570 $Y=105840
X1297 1 2 573 35 ICV_21 $T=295780 116960 0 0 $X=295590 $Y=116720
X1298 1 2 583 12 ICV_21 $T=309120 100640 0 0 $X=308930 $Y=100400
X1299 1 2 584 12 ICV_21 $T=309120 116960 0 0 $X=308930 $Y=116720
X1300 1 2 571 269 ICV_21 $T=318320 84320 1 0 $X=318130 $Y=81360
X1301 1 2 273 12 ICV_21 $T=328900 122400 1 0 $X=328710 $Y=119440
X1302 1 2 11 12 ICV_21 $T=333040 122400 0 0 $X=332850 $Y=122160
X1303 1 2 12 ICV_22 $T=6900 122400 0 0 $X=6710 $Y=122160
X1304 1 2 406 ICV_22 $T=8740 122400 1 0 $X=8550 $Y=119440
X1305 1 2 17 ICV_22 $T=12420 95200 0 0 $X=12230 $Y=94960
X1306 1 2 410 ICV_22 $T=14260 100640 1 0 $X=14070 $Y=97680
X1307 1 2 17 ICV_22 $T=17940 111520 0 0 $X=17750 $Y=111280
X1308 1 2 34 ICV_22 $T=34040 116960 0 0 $X=33850 $Y=116720
X1309 1 2 428 ICV_22 $T=34960 111520 1 0 $X=34770 $Y=108560
X1310 1 2 37 ICV_22 $T=35880 106080 0 0 $X=35690 $Y=105840
X1311 1 2 41 ICV_22 $T=38180 84320 1 0 $X=37990 $Y=81360
X1312 1 2 71 ICV_22 $T=78200 122400 0 0 $X=78010 $Y=122160
X1313 1 2 463 ICV_22 $T=100280 89760 0 0 $X=100090 $Y=89520
X1314 1 2 476 ICV_22 $T=114540 106080 0 0 $X=114350 $Y=105840
X1315 1 2 12 ICV_22 $T=118220 116960 0 0 $X=118030 $Y=116720
X1316 1 2 84 ICV_22 $T=123740 122400 1 0 $X=123550 $Y=119440
X1317 1 2 110 ICV_22 $T=131100 111520 0 0 $X=130910 $Y=111280
X1318 1 2 502 ICV_22 $T=142600 84320 0 0 $X=142410 $Y=84080
X1319 1 2 503 ICV_22 $T=142600 111520 0 0 $X=142410 $Y=111280
X1320 1 2 503 ICV_22 $T=148120 111520 0 0 $X=147930 $Y=111280
X1321 1 2 512 ICV_22 $T=163760 78880 0 0 $X=163570 $Y=78640
X1322 1 2 158 ICV_22 $T=181700 116960 0 0 $X=181510 $Y=116720
X1323 1 2 158 ICV_22 $T=211600 116960 0 0 $X=211410 $Y=116720
X1324 1 2 192 ICV_22 $T=226780 78880 0 0 $X=226590 $Y=78640
X1325 1 2 193 ICV_22 $T=226780 122400 0 0 $X=226590 $Y=122160
X1326 1 2 189 ICV_22 $T=234140 122400 0 0 $X=233950 $Y=122160
X1327 1 2 213 ICV_22 $T=246560 84320 1 0 $X=246370 $Y=81360
X1328 1 2 12 ICV_22 $T=254840 111520 0 0 $X=254650 $Y=111280
X1329 1 2 232 ICV_22 $T=269100 84320 1 0 $X=268910 $Y=81360
X1330 1 2 560 ICV_22 $T=269100 122400 1 0 $X=268910 $Y=119440
X1331 1 2 179 ICV_22 $T=273700 111520 0 0 $X=273510 $Y=111280
X1332 1 2 35 ICV_22 $T=300840 111520 1 0 $X=300650 $Y=108560
X1333 1 2 40 ICV_22 $T=302680 106080 1 0 $X=302490 $Y=103120
X1334 1 2 587 ICV_22 $T=318320 111520 1 0 $X=318130 $Y=108560
X1335 1 2 ICV_23 $T=6900 111520 0 0 $X=6710 $Y=111280
X1336 1 2 ICV_23 $T=53360 122400 1 0 $X=53170 $Y=119440
X1337 1 2 ICV_23 $T=56120 89760 1 0 $X=55930 $Y=86800
X1338 1 2 ICV_23 $T=67160 95200 0 0 $X=66970 $Y=94960
X1339 1 2 ICV_23 $T=80040 116960 1 0 $X=79850 $Y=114000
X1340 1 2 ICV_23 $T=104420 100640 1 0 $X=104230 $Y=97680
X1341 1 2 ICV_23 $T=137540 111520 1 0 $X=137350 $Y=108560
X1342 1 2 ICV_23 $T=138460 106080 1 0 $X=138270 $Y=103120
X1343 1 2 ICV_23 $T=147660 116960 1 0 $X=147470 $Y=114000
X1344 1 2 ICV_23 $T=148580 111520 1 0 $X=148390 $Y=108560
X1345 1 2 ICV_23 $T=162840 106080 1 0 $X=162650 $Y=103120
X1346 1 2 ICV_23 $T=165600 116960 1 0 $X=165410 $Y=114000
X1347 1 2 ICV_23 $T=166060 111520 1 0 $X=165870 $Y=108560
X1348 1 2 ICV_23 $T=174340 111520 0 0 $X=174150 $Y=111280
X1349 1 2 ICV_23 $T=176640 116960 1 0 $X=176450 $Y=114000
X1350 1 2 ICV_23 $T=188600 106080 1 0 $X=188410 $Y=103120
X1351 1 2 ICV_23 $T=205160 95200 1 0 $X=204970 $Y=92240
X1352 1 2 ICV_23 $T=212060 78880 0 0 $X=211870 $Y=78640
X1353 1 2 ICV_23 $T=216660 84320 1 0 $X=216470 $Y=81360
X1354 1 2 ICV_23 $T=216660 84320 0 0 $X=216470 $Y=84080
X1355 1 2 ICV_23 $T=216660 89760 1 0 $X=216470 $Y=86800
X1356 1 2 ICV_23 $T=216660 116960 1 0 $X=216470 $Y=114000
X1357 1 2 ICV_23 $T=230460 100640 0 0 $X=230270 $Y=100400
X1358 1 2 ICV_23 $T=241500 100640 0 0 $X=241310 $Y=100400
X1359 1 2 ICV_23 $T=244720 106080 1 0 $X=244530 $Y=103120
X1360 1 2 ICV_23 $T=247020 111520 1 0 $X=246830 $Y=108560
X1361 1 2 ICV_23 $T=258520 106080 0 0 $X=258330 $Y=105840
X1362 1 2 ICV_23 $T=261280 111520 1 0 $X=261090 $Y=108560
X1363 1 2 ICV_23 $T=270020 100640 0 0 $X=269830 $Y=100400
X1364 1 2 ICV_23 $T=272780 106080 1 0 $X=272590 $Y=103120
X1365 1 2 ICV_23 $T=279680 116960 1 0 $X=279490 $Y=114000
X1366 1 2 ICV_23 $T=283820 106080 1 0 $X=283630 $Y=103120
X1367 1 2 ICV_23 $T=286580 106080 0 0 $X=286390 $Y=105840
X1368 1 2 ICV_23 $T=299920 95200 0 0 $X=299730 $Y=94960
X1369 1 2 ICV_23 $T=300840 95200 1 0 $X=300650 $Y=92240
X1370 1 2 ICV_23 $T=300840 100640 1 0 $X=300650 $Y=97680
X1371 1 2 ICV_23 $T=311880 95200 1 0 $X=311690 $Y=92240
X1372 1 2 ICV_23 $T=314640 111520 0 0 $X=314450 $Y=111280
X1373 1 2 ICV_24 $T=46460 89760 1 0 $X=46270 $Y=86800
X1374 1 2 ICV_24 $T=46460 111520 1 0 $X=46270 $Y=108560
X1375 1 2 ICV_24 $T=60260 84320 0 0 $X=60070 $Y=84080
X1376 1 2 ICV_24 $T=60260 116960 0 0 $X=60070 $Y=116720
X1377 1 2 ICV_24 $T=74520 84320 1 0 $X=74330 $Y=81360
X1378 1 2 ICV_24 $T=88320 116960 0 0 $X=88130 $Y=116720
X1379 1 2 ICV_24 $T=116380 122400 0 0 $X=116190 $Y=122160
X1380 1 2 ICV_24 $T=130640 100640 1 0 $X=130450 $Y=97680
X1381 1 2 ICV_24 $T=158700 89760 1 0 $X=158510 $Y=86800
X1382 1 2 ICV_24 $T=158700 106080 1 0 $X=158510 $Y=103120
X1383 1 2 ICV_24 $T=158700 116960 1 0 $X=158510 $Y=114000
X1384 1 2 ICV_24 $T=172500 100640 0 0 $X=172310 $Y=100400
X1385 1 2 ICV_24 $T=186760 84320 1 0 $X=186570 $Y=81360
X1386 1 2 ICV_24 $T=186760 89760 1 0 $X=186570 $Y=86800
X1387 1 2 ICV_24 $T=228620 89760 0 0 $X=228430 $Y=89520
X1388 1 2 ICV_24 $T=242880 106080 1 0 $X=242690 $Y=103120
X1389 1 2 ICV_24 $T=256680 106080 0 0 $X=256490 $Y=105840
X1390 1 2 ICV_24 $T=299000 89760 1 0 $X=298810 $Y=86800
X1391 1 2 ICV_24 $T=312800 122400 0 0 $X=312610 $Y=122160
X1392 1 2 ICV_24 $T=327060 100640 1 0 $X=326870 $Y=97680
X1393 1 2 ICV_24 $T=327060 116960 1 0 $X=326870 $Y=114000
X1394 1 2 ICV_29 $T=10580 106080 1 0 $X=10390 $Y=103120
X1395 1 2 ICV_29 $T=10580 111520 1 0 $X=10390 $Y=108560
X1396 1 2 ICV_29 $T=10580 116960 1 0 $X=10390 $Y=114000
X1397 1 2 ICV_29 $T=18400 106080 0 0 $X=18210 $Y=105840
X1398 1 2 ICV_29 $T=37260 111520 1 0 $X=37070 $Y=108560
X1399 1 2 ICV_29 $T=38640 95200 1 0 $X=38450 $Y=92240
X1400 1 2 ICV_29 $T=53820 106080 1 0 $X=53630 $Y=103120
X1401 1 2 ICV_29 $T=67160 84320 0 0 $X=66970 $Y=84080
X1402 1 2 ICV_29 $T=79120 116960 0 0 $X=78930 $Y=116720
X1403 1 2 ICV_29 $T=114540 122400 1 0 $X=114350 $Y=119440
X1404 1 2 ICV_29 $T=121900 111520 0 0 $X=121710 $Y=111280
X1405 1 2 ICV_29 $T=126040 106080 0 0 $X=125850 $Y=105840
X1406 1 2 ICV_29 $T=133400 111520 0 0 $X=133210 $Y=111280
X1407 1 2 ICV_29 $T=149500 106080 1 0 $X=149310 $Y=103120
X1408 1 2 ICV_29 $T=188600 100640 0 0 $X=188410 $Y=100400
X1409 1 2 ICV_29 $T=206540 100640 1 0 $X=206350 $Y=97680
X1410 1 2 ICV_29 $T=219420 89760 0 0 $X=219230 $Y=89520
X1411 1 2 ICV_29 $T=269560 106080 0 0 $X=269370 $Y=105840
X1412 1 2 ICV_29 $T=303600 122400 0 0 $X=303410 $Y=122160
X1413 1 2 ICV_29 $T=323840 95200 0 0 $X=323650 $Y=94960
X1414 1 2 438 430 2 28 1 sky130_fd_sc_hd__or2_4 $T=46920 106080 0 0 $X=46730 $Y=105840
X1415 1 2 438 43 2 31 1 sky130_fd_sc_hd__or2_4 $T=49220 89760 1 0 $X=49030 $Y=86800
X1416 1 2 438 47 2 49 1 sky130_fd_sc_hd__or2_4 $T=50600 106080 1 0 $X=50410 $Y=103120
X1417 1 2 438 48 2 34 1 sky130_fd_sc_hd__or2_4 $T=51060 100640 0 0 $X=50870 $Y=100400
X1418 1 2 438 44 2 33 1 sky130_fd_sc_hd__or2_4 $T=52440 95200 0 0 $X=52250 $Y=94960
X1419 1 2 50 429 2 39 1 sky130_fd_sc_hd__or2_4 $T=54280 106080 0 0 $X=54090 $Y=105840
X1420 1 2 50 62 2 63 1 sky130_fd_sc_hd__or2_4 $T=65780 122400 1 0 $X=65590 $Y=119440
X1421 1 2 73 61 2 74 1 sky130_fd_sc_hd__or2_4 $T=84640 89760 1 0 $X=84450 $Y=86800
X1422 1 2 463 468 2 446 1 sky130_fd_sc_hd__or2_4 $T=89240 95200 1 0 $X=89050 $Y=92240
X1423 1 2 458 468 2 64 1 sky130_fd_sc_hd__or2_4 $T=91080 89760 0 0 $X=90890 $Y=89520
X1424 1 2 464 468 2 450 1 sky130_fd_sc_hd__or2_4 $T=91080 100640 0 0 $X=90890 $Y=100400
X1425 1 2 466 468 2 461 1 sky130_fd_sc_hd__or2_4 $T=92000 106080 0 0 $X=91810 $Y=105840
X1426 1 2 75 76 2 81 1 sky130_fd_sc_hd__or2_4 $T=93840 116960 1 0 $X=93650 $Y=114000
X1427 1 2 467 468 2 462 1 sky130_fd_sc_hd__or2_4 $T=94300 100640 1 0 $X=94110 $Y=97680
X1428 1 2 472 90 2 465 1 sky130_fd_sc_hd__or2_4 $T=109940 95200 0 0 $X=109750 $Y=94960
X1429 1 2 89 90 2 97 1 sky130_fd_sc_hd__or2_4 $T=110860 84320 0 0 $X=110670 $Y=84080
X1430 1 2 105 479 2 106 1 sky130_fd_sc_hd__or2_4 $T=124660 122400 0 0 $X=124470 $Y=122160
X1431 1 2 105 99 2 116 1 sky130_fd_sc_hd__or2_4 $T=135700 116960 0 0 $X=135510 $Y=116720
X1432 1 2 503 491 2 120 1 sky130_fd_sc_hd__or2_4 $T=144440 116960 1 0 $X=144250 $Y=114000
X1433 1 2 503 127 2 129 1 sky130_fd_sc_hd__or2_4 $T=151340 111520 0 0 $X=151150 $Y=111280
X1434 1 2 503 132 2 133 1 sky130_fd_sc_hd__or2_4 $T=154100 106080 0 0 $X=153910 $Y=105840
X1435 1 2 503 139 2 143 1 sky130_fd_sc_hd__or2_4 $T=162380 116960 1 0 $X=162190 $Y=114000
X1436 1 2 518 156 2 511 1 sky130_fd_sc_hd__or2_4 $T=179400 95200 1 0 $X=179210 $Y=92240
X1437 1 2 155 108 2 512 1 sky130_fd_sc_hd__or2_4 $T=179860 84320 1 0 $X=179670 $Y=81360
X1438 1 2 520 151 2 513 1 sky130_fd_sc_hd__or2_4 $T=179860 89760 1 0 $X=179670 $Y=86800
X1439 1 2 87 160 2 388 1 sky130_fd_sc_hd__or2_4 $T=183540 89760 0 0 $X=183350 $Y=89520
X1440 1 2 9 152 2 389 1 sky130_fd_sc_hd__or2_4 $T=202400 84320 1 0 $X=202210 $Y=81360
X1441 1 2 522 172 2 525 1 sky130_fd_sc_hd__or2_4 $T=202860 89760 1 0 $X=202670 $Y=86800
X1442 1 2 180 160 2 518 1 sky130_fd_sc_hd__or2_4 $T=209300 84320 1 0 $X=209110 $Y=81360
X1443 1 2 244 191 2 251 1 sky130_fd_sc_hd__or2_4 $T=294400 78880 0 0 $X=294210 $Y=78640
X1444 1 2 240 527 2 256 1 sky130_fd_sc_hd__or2_4 $T=301760 89760 1 0 $X=301570 $Y=86800
X1445 1 2 242 527 2 582 1 sky130_fd_sc_hd__or2_4 $T=303600 89760 0 0 $X=303410 $Y=89520
X1446 1 2 498 397 2 517 1 sky130_fd_sc_hd__and2_4 $T=172960 89760 1 0 $X=172770 $Y=86800
X1447 1 2 122 159 2 6 1 sky130_fd_sc_hd__and2_4 $T=189060 84320 0 0 $X=188870 $Y=84080
X1448 1 2 5 523 2 524 1 sky130_fd_sc_hd__and2_4 $T=195960 89760 1 0 $X=195770 $Y=86800
X1449 1 2 7 161 2 527 1 sky130_fd_sc_hd__and2_4 $T=199640 100640 1 0 $X=199450 $Y=97680
X1450 1 2 221 216 2 543 1 sky130_fd_sc_hd__and2_4 $T=256220 89760 1 0 $X=256030 $Y=86800
X1451 1 2 224 230 2 211 1 sky130_fd_sc_hd__and2_4 $T=266340 78880 0 0 $X=266150 $Y=78640
X1452 1 2 258 544 2 579 1 sky130_fd_sc_hd__and2_4 $T=306820 84320 0 0 $X=306630 $Y=84080
X1453 1 2 269 571 2 270 1 sky130_fd_sc_hd__and2_4 $T=319700 89760 1 0 $X=319510 $Y=86800
X1454 1 2 176 524 515 2 530 1 sky130_fd_sc_hd__nor3_4 $T=203320 84320 0 0 $X=203130 $Y=84080
X1455 1 2 215 547 550 2 551 1 sky130_fd_sc_hd__nor3_4 $T=252080 100640 1 0 $X=251890 $Y=97680
X1456 1 2 255 579 257 2 260 1 sky130_fd_sc_hd__nor3_4 $T=303600 78880 0 0 $X=303410 $Y=78640
X1457 1 2 255 270 263 2 265 1 sky130_fd_sc_hd__nor3_4 $T=315560 78880 0 0 $X=315370 $Y=78640
X1458 1 2 6 145 113 164 2 1 sky130_fd_sc_hd__a21oi_4 $T=192280 78880 0 0 $X=192090 $Y=78640
X1459 1 2 228 555 559 558 2 1 sky130_fd_sc_hd__a21oi_4 $T=265420 95200 0 0 $X=265230 $Y=94960
X1460 1 2 582 267 261 263 2 1 sky130_fd_sc_hd__a21oi_4 $T=312340 84320 1 0 $X=312150 $Y=81360
X1461 1 12 425 ICV_36 $T=29900 100640 0 0 $X=29710 $Y=100400
X1462 1 51 41 ICV_36 $T=57960 111520 0 0 $X=57770 $Y=111280
X1463 1 463 458 ICV_36 $T=86020 89760 0 0 $X=85830 $Y=89520
X1464 1 460 460 ICV_36 $T=86020 95200 0 0 $X=85830 $Y=94960
X1465 1 460 468 ICV_36 $T=86020 100640 0 0 $X=85830 $Y=100400
X1466 1 90 491 ICV_36 $T=114080 95200 0 0 $X=113890 $Y=94960
X1467 1 508 506 ICV_36 $T=156400 95200 1 0 $X=156210 $Y=92240
X1468 1 513 148 ICV_36 $T=170200 89760 0 0 $X=170010 $Y=89520
X1469 1 514 12 ICV_36 $T=170200 122400 0 0 $X=170010 $Y=122160
X1470 1 172 522 ICV_36 $T=198260 84320 0 0 $X=198070 $Y=84080
X1471 1 7 392 ICV_36 $T=198260 100640 0 0 $X=198070 $Y=100400
X1472 1 166 175 ICV_36 $T=198260 111520 0 0 $X=198070 $Y=111280
X1473 1 548 222 ICV_36 $T=254380 78880 0 0 $X=254190 $Y=78640
X1474 1 201 216 ICV_36 $T=254380 84320 0 0 $X=254190 $Y=84080
X1475 1 559 220 ICV_36 $T=268640 89760 1 0 $X=268450 $Y=86800
X1476 1 261 255 ICV_36 $T=310500 78880 0 0 $X=310310 $Y=78640
X1477 1 167 578 ICV_36 $T=310500 111520 0 0 $X=310310 $Y=111280
X1478 1 2 65 67 65 439 ICV_37 $T=69920 78880 0 0 $X=69730 $Y=78640
X1479 1 2 87 90 87 468 ICV_37 $T=104880 84320 0 0 $X=104690 $Y=84080
X1480 1 2 128 508 508 113 ICV_37 $T=158700 78880 0 0 $X=158510 $Y=78640
X1481 1 2 131 507 507 500 ICV_37 $T=159620 95200 0 0 $X=159430 $Y=94960
X1482 1 2 459 12 459 146 ICV_37 $T=166060 95200 0 0 $X=165870 $Y=94960
X1483 1 2 511 511 511 459 ICV_37 $T=166060 106080 0 0 $X=165870 $Y=105840
X1484 1 2 130 114 130 122 ICV_37 $T=166980 78880 0 0 $X=166790 $Y=78640
X1485 1 2 519 163 519 162 ICV_37 $T=188600 122400 0 0 $X=188410 $Y=122160
X1486 1 2 161 519 519 3 ICV_37 $T=189520 106080 0 0 $X=189330 $Y=105840
X1487 1 2 12 30 30 167 ICV_37 $T=194580 122400 0 0 $X=194390 $Y=122160
X1488 1 2 392 433 433 177 ICV_37 $T=203780 116960 1 0 $X=203590 $Y=114000
X1489 1 2 538 197 538 36 ICV_37 $T=231380 111520 0 0 $X=231190 $Y=111280
X1490 1 2 206 518 518 537 ICV_37 $T=234600 89760 0 0 $X=234410 $Y=89520
X1491 1 2 232 232 548 559 ICV_37 $T=273700 89760 1 0 $X=273510 $Y=86800
X1492 1 2 546 546 567 199 ICV_37 $T=292100 95200 1 0 $X=291910 $Y=92240
X1493 1 2 568 567 568 248 ICV_37 $T=294400 89760 0 0 $X=294210 $Y=89520
X1494 1 2 579 257 527 244 ICV_37 $T=301760 84320 1 0 $X=301570 $Y=81360
X1495 1 2 497 112 499 500 2 467 1 sky130_fd_sc_hd__or4_4 $T=135700 100640 0 0 $X=135510 $Y=100400
X1496 1 2 497 112 501 500 2 472 1 sky130_fd_sc_hd__or4_4 $T=136160 89760 0 0 $X=135970 $Y=89520
X1497 1 2 497 111 499 502 2 463 1 sky130_fd_sc_hd__or4_4 $T=136160 95200 0 0 $X=135970 $Y=94960
X1498 1 2 114 112 499 500 2 117 1 sky130_fd_sc_hd__or4_4 $T=136620 84320 0 0 $X=136430 $Y=84080
X1499 1 2 497 111 501 502 2 466 1 sky130_fd_sc_hd__or4_4 $T=137080 100640 1 0 $X=136890 $Y=97680
X1500 1 2 113 498 107 115 2 118 1 sky130_fd_sc_hd__or4_4 $T=138000 78880 0 0 $X=137810 $Y=78640
X1501 1 2 107 115 499 502 2 89 1 sky130_fd_sc_hd__or4_4 $T=138460 95200 1 0 $X=138270 $Y=92240
X1502 1 2 108 114 501 498 2 119 1 sky130_fd_sc_hd__or4_4 $T=139380 84320 1 0 $X=139190 $Y=81360
X1503 1 2 108 504 499 109 2 458 1 sky130_fd_sc_hd__or4_4 $T=139840 89760 1 0 $X=139650 $Y=86800
X1504 1 2 107 504 501 500 2 505 1 sky130_fd_sc_hd__or4_4 $T=146280 95200 1 0 $X=146090 $Y=92240
X1505 1 2 108 114 122 498 2 123 1 sky130_fd_sc_hd__or4_4 $T=147200 78880 0 0 $X=147010 $Y=78640
X1506 1 2 122 109 107 115 2 124 1 sky130_fd_sc_hd__or4_4 $T=147200 84320 1 0 $X=147010 $Y=81360
X1507 1 2 504 112 501 502 2 125 1 sky130_fd_sc_hd__or4_4 $T=147200 89760 0 0 $X=147010 $Y=89520
X1508 1 2 506 115 508 507 2 137 1 sky130_fd_sc_hd__or4_4 $T=155480 89760 0 0 $X=155290 $Y=89520
X1509 1 2 504 128 130 131 2 136 1 sky130_fd_sc_hd__or4_4 $T=155940 84320 0 0 $X=155750 $Y=84080
X1510 1 2 519 152 113 109 2 155 1 sky130_fd_sc_hd__or4_4 $T=181240 84320 0 0 $X=181050 $Y=84080
X1511 1 2 543 214 213 211 2 521 1 sky130_fd_sc_hd__or4_4 $T=245640 84320 0 0 $X=245450 $Y=84080
X1512 1 2 201 214 213 211 2 544 1 sky130_fd_sc_hd__or4_4 $T=259440 84320 0 0 $X=259250 $Y=84080
X1513 1 2 219 220 546 9 2 556 1 sky130_fd_sc_hd__or4_4 $T=259440 89760 0 0 $X=259250 $Y=89520
X1514 1 2 221 222 227 172 2 557 1 sky130_fd_sc_hd__or4_4 $T=263120 84320 1 0 $X=262930 $Y=81360
X1515 1 2 235 559 232 233 2 566 1 sky130_fd_sc_hd__or4_4 $T=277840 84320 0 0 $X=277650 $Y=84080
X1516 1 2 235 559 221 564 2 567 1 sky130_fd_sc_hd__or4_4 $T=278300 89760 0 0 $X=278110 $Y=89520
X1517 1 2 235 559 232 220 2 568 1 sky130_fd_sc_hd__or4_4 $T=279680 89760 1 0 $X=279490 $Y=86800
X1518 1 2 235 559 221 233 2 569 1 sky130_fd_sc_hd__or4_4 $T=287500 89760 0 0 $X=287310 $Y=89520
X1519 1 2 498 122 108 2 154 1 sky130_fd_sc_hd__and3_4 $T=175260 78880 0 0 $X=175070 $Y=78640
X1520 1 2 224 548 222 2 216 1 sky130_fd_sc_hd__and3_4 $T=259440 78880 0 0 $X=259250 $Y=78640
X1521 1 2 233 232 230 2 209 1 sky130_fd_sc_hd__and3_4 $T=273240 78880 0 0 $X=273050 $Y=78640
X1522 1 2 233 219 230 2 237 1 sky130_fd_sc_hd__and3_4 $T=281060 84320 1 0 $X=280870 $Y=81360
X1523 1 2 220 232 230 2 570 1 sky130_fd_sc_hd__and3_4 $T=287500 78880 0 0 $X=287310 $Y=78640
X1524 1 2 497 8 168 2 523 1 sky130_fd_sc_hd__or3_4 $T=203320 95200 0 0 $X=203130 $Y=94960
X1525 1 2 216 213 211 2 206 1 sky130_fd_sc_hd__or3_4 $T=248400 89760 1 0 $X=248210 $Y=86800
X1526 1 2 214 211 216 2 207 1 sky130_fd_sc_hd__or3_4 $T=249780 84320 1 0 $X=249590 $Y=81360
X1527 1 2 122 159 109 93 2 520 1 sky130_fd_sc_hd__and4_4 $T=183080 78880 0 0 $X=182890 $Y=78640
X1528 1 2 142 512 114 2 515 1 sky130_fd_sc_hd__a21boi_4 $T=169280 84320 1 0 $X=169090 $Y=81360
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_1 VNB VPB A X VPWR VGND
** N=18 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 VGND 7 X VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=395 $Y=235 $D=9
M1 7 A VGND VNB nshort L=0.15 W=0.52 m=1 r=3.46667 a=0.078 p=1.34 mult=1 $X=835 $Y=235 $D=9
M2 VPWR 7 X VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=395 $Y=1695 $D=89
M3 7 A VPWR VPB phighvt L=0.15 W=0.79 m=1 r=5.26667 a=0.1185 p=1.88 mult=1 $X=835 $Y=1695 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_4 VNB VPB A VPWR X VGND
** N=28 EP=6 IP=0 FDC=10
*.SEEDPROM
M0 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=885 $Y=235 $D=9
M2 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1315 $Y=235 $D=9
M3 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1745 $Y=235 $D=9
M4 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2175 $Y=235 $D=9
M5 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M6 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=880 $Y=1485 $D=89
M7 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1310 $Y=1485 $D=89
M8 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M9 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_16 VNB VPB A VPWR X VGND
** N=79 EP=6 IP=0 FDC=40
*.SEEDPROM
M0 7 A VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=830 $Y=235 $D=9
M2 7 A VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1260 $Y=235 $D=9
M3 VGND A 7 VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=1690 $Y=235 $D=9
M4 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2120 $Y=235 $D=9
M5 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2550 $Y=235 $D=9
M6 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=2980 $Y=235 $D=9
M7 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3410 $Y=235 $D=9
M8 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=3840 $Y=235 $D=9
M9 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4270 $Y=235 $D=9
M10 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=4700 $Y=235 $D=9
M11 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5130 $Y=235 $D=9
M12 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5555 $Y=235 $D=9
M13 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=5985 $Y=235 $D=9
M14 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M15 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=6845 $Y=235 $D=9
M16 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7275 $Y=235 $D=9
M17 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=7705 $Y=235 $D=9
M18 X 7 VGND VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8135 $Y=235 $D=9
M19 VGND 7 X VNB nshort L=0.15 W=0.42 m=1 r=2.8 a=0.063 p=1.14 mult=1 $X=8565 $Y=235 $D=9
M20 7 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M21 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M22 7 A VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M23 VPWR A 7 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M24 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2120 $Y=1485 $D=89
M25 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2550 $Y=1485 $D=89
M26 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2980 $Y=1485 $D=89
M27 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3410 $Y=1485 $D=89
M28 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3840 $Y=1485 $D=89
M29 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4270 $Y=1485 $D=89
M30 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4700 $Y=1485 $D=89
M31 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5130 $Y=1485 $D=89
M32 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5555 $Y=1485 $D=89
M33 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=5985 $Y=1485 $D=89
M34 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6415 $Y=1485 $D=89
M35 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6845 $Y=1485 $D=89
M36 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
M37 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7705 $Y=1485 $D=89
M38 X 7 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8135 $Y=1485 $D=89
M39 VPWR 7 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=8565 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a21o_4 VNB VPB B1 A2 A1 VPWR X VGND
** N=55 EP=8 IP=0 FDC=20
*.SEEDPROM
M0 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=420 $Y=235 $D=9
M1 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=850 $Y=235 $D=9
M2 X 9 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1280 $Y=235 $D=9
M3 VGND 9 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1710 $Y=235 $D=9
M4 9 B1 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2675 $Y=235 $D=9
M5 VGND B1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3095 $Y=235 $D=9
M6 11 A2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3555 $Y=235 $D=9
M7 9 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3935 $Y=235 $D=9
M8 12 A1 9 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4355 $Y=235 $D=9
M9 VGND A2 12 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4775 $Y=235 $D=9
M10 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=420 $Y=1485 $D=89
M11 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=850 $Y=1485 $D=89
M12 X 9 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1280 $Y=1485 $D=89
M13 VPWR 9 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1710 $Y=1485 $D=89
M14 9 B1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2675 $Y=1485 $D=89
M15 10 B1 9 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3095 $Y=1485 $D=89
M16 VPWR A2 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3515 $Y=1485 $D=89
M17 10 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3935 $Y=1485 $D=89
M18 VPWR A1 10 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4355 $Y=1485 $D=89
M19 10 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4775 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4
** N=4 EP=4 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=2760 0 0 0 $X=2570 $Y=-240
X1 1 3 4 ICV_7 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__a32o_4 VNB VPB A3 A2 A1 B1 B2 VPWR X VGND
** N=67 EP=10 IP=0 FDC=28
*.SEEDPROM
M0 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 X 11 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 VGND 11 X VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 13 A3 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2075 $Y=235 $D=9
M5 VGND A3 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=2495 $Y=235 $D=9
M6 13 A2 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3435 $Y=235 $D=9
M7 14 A2 13 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=3855 $Y=235 $D=9
M8 11 A1 14 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4275 $Y=235 $D=9
M9 14 A1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=4695 $Y=235 $D=9
M10 11 B1 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=5970 $Y=235 $D=9
M11 15 B1 11 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6390 $Y=235 $D=9
M12 VGND B2 15 VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=6855 $Y=235 $D=9
M13 15 B2 VGND VNB nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=7275 $Y=235 $D=9
M14 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M15 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M16 X 11 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M17 VPWR 11 X VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M18 12 A3 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2075 $Y=1485 $D=89
M19 VPWR A3 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=2495 $Y=1485 $D=89
M20 VPWR A2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3435 $Y=1485 $D=89
M21 12 A2 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=3855 $Y=1485 $D=89
M22 VPWR A1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4275 $Y=1485 $D=89
M23 12 A1 VPWR VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=4695 $Y=1485 $D=89
M24 11 B1 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6015 $Y=1485 $D=89
M25 12 B1 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6435 $Y=1485 $D=89
M26 11 B2 12 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=6855 $Y=1485 $D=89
M27 12 B2 11 VPB phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257
** N=733 EP=257 IP=5958 FDC=8220
M0 1 328 339 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=183015 $Y=57355 $D=9
M1 339 328 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=183435 $Y=57355 $D=9
M2 1 328 339 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=183855 $Y=57355 $D=9
M3 339 328 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=184275 $Y=57355 $D=9
M4 334 3 339 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=184695 $Y=57355 $D=9
M5 339 3 334 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=185115 $Y=57355 $D=9
M6 334 3 339 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=185535 $Y=57355 $D=9
M7 339 3 334 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=185955 $Y=57355 $D=9
M8 334 329 340 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=186895 $Y=57355 $D=9
M9 340 329 334 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=187315 $Y=57355 $D=9
M10 334 329 340 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=187735 $Y=57355 $D=9
M11 340 329 334 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=188155 $Y=57355 $D=9
M12 341 330 340 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=188715 $Y=57355 $D=9
M13 340 330 341 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=189135 $Y=57355 $D=9
M14 341 330 340 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=189555 $Y=57355 $D=9
M15 340 330 341 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=189975 $Y=57355 $D=9
M16 341 4 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=190915 $Y=57355 $D=9
M17 1 4 341 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=191335 $Y=57355 $D=9
M18 341 4 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=191755 $Y=57355 $D=9
M19 1 4 341 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=192175 $Y=57355 $D=9
M20 338 5 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=203735 $Y=68235 $D=9
M21 1 5 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204155 $Y=68235 $D=9
M22 338 5 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204575 $Y=68235 $D=9
M23 1 5 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=204995 $Y=68235 $D=9
M24 338 6 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=205415 $Y=68235 $D=9
M25 1 6 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=205835 $Y=68235 $D=9
M26 338 6 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=206255 $Y=68235 $D=9
M27 1 6 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=206675 $Y=68235 $D=9
M28 338 331 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=207615 $Y=68235 $D=9
M29 1 331 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=208035 $Y=68235 $D=9
M30 338 331 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=208455 $Y=68235 $D=9
M31 1 331 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=208875 $Y=68235 $D=9
M32 338 332 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=209295 $Y=68235 $D=9
M33 1 332 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=209715 $Y=68235 $D=9
M34 338 332 1 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=210135 $Y=68235 $D=9
M35 1 332 338 1 nshort L=0.15 W=0.65 m=1 r=4.33333 a=0.0975 p=1.6 mult=1 $X=210555 $Y=68235 $D=9
M36 334 328 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=183015 $Y=58605 $D=89
M37 333 328 334 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=183435 $Y=58605 $D=89
M38 334 328 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=183855 $Y=58605 $D=89
M39 333 328 334 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=184275 $Y=58605 $D=89
M40 334 3 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=184695 $Y=58605 $D=89
M41 333 3 334 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=185115 $Y=58605 $D=89
M42 334 3 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=185535 $Y=58605 $D=89
M43 333 3 334 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=185955 $Y=58605 $D=89
M44 2 329 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=186395 $Y=58605 $D=89
M45 333 329 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=186815 $Y=58605 $D=89
M46 2 329 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=187235 $Y=58605 $D=89
M47 333 329 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=188060 $Y=58605 $D=89
M48 2 330 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=188715 $Y=58605 $D=89
M49 333 330 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=189135 $Y=58605 $D=89
M50 2 330 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=189555 $Y=58605 $D=89
M51 333 330 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=189975 $Y=58605 $D=89
M52 2 4 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=190915 $Y=58605 $D=89
M53 333 4 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=191335 $Y=58605 $D=89
M54 2 4 333 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=191755 $Y=58605 $D=89
M55 333 4 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=192175 $Y=58605 $D=89
M56 2 5 335 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=203735 $Y=69485 $D=89
M57 335 5 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204155 $Y=69485 $D=89
M58 2 5 335 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204575 $Y=69485 $D=89
M59 335 5 2 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=204995 $Y=69485 $D=89
M60 336 6 335 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=205415 $Y=69485 $D=89
M61 335 6 336 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=205835 $Y=69485 $D=89
M62 336 6 335 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=206255 $Y=69485 $D=89
M63 335 6 336 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=206675 $Y=69485 $D=89
M64 336 331 337 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=207615 $Y=69485 $D=89
M65 337 331 336 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=208035 $Y=69485 $D=89
M66 336 331 337 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=208455 $Y=69485 $D=89
M67 337 331 336 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=208875 $Y=69485 $D=89
M68 338 332 337 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=209295 $Y=69485 $D=89
M69 337 332 338 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=209715 $Y=69485 $D=89
M70 338 332 337 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=210135 $Y=69485 $D=89
M71 337 332 338 2 phighvt L=0.15 W=1 m=1 r=6.66667 a=0.15 p=2.3 mult=1 $X=210555 $Y=69485 $D=89
X72 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=36665 $D=191
X73 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=42105 $D=191
X74 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=47545 $D=191
X75 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=52985 $D=191
X76 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=58425 $D=191
X77 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=63865 $D=191
X78 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=69305 $D=191
X79 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=74745 $D=191
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 35360 0 0 $X=6710 $Y=35120
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=14260 68000 0 0 $X=14070 $Y=67760
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18860 35360 0 0 $X=18670 $Y=35120
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28520 35360 0 0 $X=28330 $Y=35120
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=31280 62560 1 0 $X=31090 $Y=59600
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=31280 73440 1 0 $X=31090 $Y=70480
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=32200 73440 0 0 $X=32010 $Y=73200
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=38640 68000 1 0 $X=38450 $Y=65040
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=42780 57120 0 0 $X=42590 $Y=56880
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=53820 51680 0 0 $X=53630 $Y=51440
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=60260 35360 0 0 $X=60070 $Y=35120
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=60260 40800 0 0 $X=60070 $Y=40560
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=60260 46240 0 0 $X=60070 $Y=46000
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=70840 57120 1 0 $X=70650 $Y=54160
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=73140 40800 0 0 $X=72950 $Y=40560
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=78660 46240 1 0 $X=78470 $Y=43280
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=86020 73440 1 0 $X=85830 $Y=70480
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88320 73440 0 0 $X=88130 $Y=73200
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=90160 68000 0 0 $X=89970 $Y=67760
X99 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=98440 51680 0 0 $X=98250 $Y=51440
X100 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 73440 1 0 $X=102390 $Y=70480
X101 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=129720 51680 0 0 $X=129530 $Y=51440
X102 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=136160 57120 1 0 $X=135970 $Y=54160
X103 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 68000 1 0 $X=158510 $Y=65040
X104 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 57120 1 0 $X=160350 $Y=54160
X105 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=172960 68000 1 0 $X=172770 $Y=65040
X106 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=181240 62560 1 0 $X=181050 $Y=59600
X107 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=197800 46240 1 0 $X=197610 $Y=43280
X108 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=197800 68000 1 0 $X=197610 $Y=65040
X109 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 40800 1 0 $X=214630 $Y=37840
X110 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 51680 1 0 $X=214630 $Y=48720
X111 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 57120 1 0 $X=214630 $Y=54160
X112 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220800 57120 0 0 $X=220610 $Y=56880
X113 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224940 40800 0 0 $X=224750 $Y=40560
X114 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224940 46240 0 0 $X=224750 $Y=46000
X115 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=226780 46240 1 0 $X=226590 $Y=43280
X116 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228620 35360 0 0 $X=228430 $Y=35120
X117 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228620 57120 0 0 $X=228430 $Y=56880
X118 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 57120 0 0 $X=230270 $Y=56880
X119 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=241040 57120 1 0 $X=240850 $Y=54160
X120 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 62560 1 0 $X=242690 $Y=59600
X121 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 73440 1 0 $X=242690 $Y=70480
X122 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=244720 57120 1 0 $X=244530 $Y=54160
X123 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=247020 51680 1 0 $X=246830 $Y=48720
X124 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 51680 1 0 $X=270750 $Y=48720
X125 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 78880 1 0 $X=270750 $Y=75920
X126 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=279220 57120 1 0 $X=279030 $Y=54160
X127 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=285200 51680 1 0 $X=285010 $Y=48720
X128 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286120 68000 1 0 $X=285930 $Y=65040
X129 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286580 68000 0 0 $X=286390 $Y=67760
X130 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 68000 1 0 $X=300650 $Y=65040
X131 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=305900 40800 0 0 $X=305710 $Y=40560
X132 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=328900 51680 1 0 $X=328710 $Y=48720
X133 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=333040 51680 0 0 $X=332850 $Y=51440
X134 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 51680 0 0 $X=340670 $Y=51440
X226 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=18400 62560 0 0 $X=18210 $Y=62320
X227 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 57120 1 0 $X=20050 $Y=54160
X228 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 68000 0 0 $X=29710 $Y=67760
X229 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=36800 73440 1 0 $X=36610 $Y=70480
X230 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39100 51680 0 0 $X=38910 $Y=51440
X231 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39100 57120 0 0 $X=38910 $Y=56880
X232 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=43700 40800 1 0 $X=43510 $Y=37840
X233 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=48300 40800 1 0 $X=48110 $Y=37840
X234 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=54280 57120 0 0 $X=54090 $Y=56880
X235 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=55660 73440 1 0 $X=55470 $Y=70480
X236 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=67160 51680 0 0 $X=66970 $Y=51440
X237 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=69460 40800 0 0 $X=69270 $Y=40560
X238 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71760 62560 0 0 $X=71570 $Y=62320
X239 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=83720 78880 1 0 $X=83530 $Y=75920
X240 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 35360 0 0 $X=89970 $Y=35120
X241 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=97520 73440 0 0 $X=97330 $Y=73200
X242 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=106260 35360 0 0 $X=106070 $Y=35120
X243 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=109940 40800 1 0 $X=109750 $Y=37840
X244 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=112240 78880 1 0 $X=112050 $Y=75920
X245 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=114540 57120 1 0 $X=114350 $Y=54160
X246 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=117300 68000 1 0 $X=117110 $Y=65040
X247 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=122360 68000 1 0 $X=122170 $Y=65040
X248 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 40800 1 0 $X=128150 $Y=37840
X249 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142600 40800 1 0 $X=142410 $Y=37840
X250 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=149040 46240 1 0 $X=148850 $Y=43280
X251 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=154100 62560 1 0 $X=153910 $Y=59600
X252 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 73440 1 0 $X=156210 $Y=70480
X253 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=164680 46240 1 0 $X=164490 $Y=43280
X254 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=177560 62560 1 0 $X=177370 $Y=59600
X255 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183540 51680 1 0 $X=183350 $Y=48720
X256 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=191360 40800 0 0 $X=191170 $Y=40560
X257 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194120 46240 1 0 $X=193930 $Y=43280
X258 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=195040 40800 1 0 $X=194850 $Y=37840
X259 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=208840 51680 0 0 $X=208650 $Y=51440
X260 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 57120 1 0 $X=210950 $Y=54160
X261 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 46240 1 0 $X=216470 $Y=43280
X262 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=224940 35360 0 0 $X=224750 $Y=35120
X263 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=237360 57120 1 0 $X=237170 $Y=54160
X264 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=244720 46240 1 0 $X=244530 $Y=43280
X265 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249320 57120 1 0 $X=249130 $Y=54160
X266 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268180 68000 1 0 $X=267990 $Y=65040
X267 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 73440 1 0 $X=268450 $Y=70480
X268 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 62560 1 0 $X=272590 $Y=59600
X269 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=276000 51680 0 0 $X=275810 $Y=51440
X270 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=277840 73440 1 0 $X=277650 $Y=70480
X271 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282440 68000 1 0 $X=282250 $Y=65040
X272 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=283360 73440 1 0 $X=283170 $Y=70480
X273 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=293480 62560 0 0 $X=293290 $Y=62320
X274 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=320160 57120 0 0 $X=319970 $Y=56880
X275 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 57120 1 0 $X=324570 $Y=54160
X276 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 78880 1 0 $X=324570 $Y=75920
X277 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 40800 1 0 $X=344810 $Y=37840
X278 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 57120 1 0 $X=344810 $Y=54160
X279 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 73440 1 0 $X=344810 $Y=70480
X280 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 46240 1 0 $X=345270 $Y=43280
X281 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 51680 1 0 $X=345270 $Y=48720
X282 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 62560 1 0 $X=345270 $Y=59600
X283 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 78880 1 0 $X=345270 $Y=75920
X284 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=14260 68000 1 0 $X=14070 $Y=65040
X285 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=18400 40800 0 0 $X=18210 $Y=40560
X286 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=18400 51680 0 0 $X=18210 $Y=51440
X287 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25300 62560 0 0 $X=25110 $Y=62320
X288 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25760 62560 1 0 $X=25570 $Y=59600
X289 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25760 73440 1 0 $X=25570 $Y=70480
X290 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=34960 57120 1 0 $X=34770 $Y=54160
X291 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=36800 62560 1 0 $X=36610 $Y=59600
X292 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40480 51680 1 0 $X=40290 $Y=48720
X293 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=40480 57120 1 0 $X=40290 $Y=54160
X294 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=41400 73440 0 0 $X=41210 $Y=73200
X295 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=42320 62560 1 0 $X=42130 $Y=59600
X296 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=45540 46240 0 0 $X=45350 $Y=46000
X297 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=51980 62560 1 0 $X=51790 $Y=59600
X298 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55660 73440 0 0 $X=55470 $Y=73200
X299 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=62560 40800 1 0 $X=62370 $Y=37840
X300 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=65780 51680 1 0 $X=65590 $Y=48720
X301 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=66700 46240 1 0 $X=66510 $Y=43280
X302 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=68080 40800 1 0 $X=67890 $Y=37840
X303 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=70380 62560 1 0 $X=70190 $Y=59600
X304 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81880 68000 1 0 $X=81690 $Y=65040
X305 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=96140 62560 1 0 $X=95950 $Y=59600
X306 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97060 73440 1 0 $X=96870 $Y=70480
X307 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97980 46240 0 0 $X=97790 $Y=46000
X308 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97980 68000 1 0 $X=97790 $Y=65040
X309 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=109480 46240 1 0 $X=109290 $Y=43280
X310 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=117300 62560 1 0 $X=117110 $Y=59600
X311 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=132020 35360 0 0 $X=131830 $Y=35120
X312 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=138460 40800 0 0 $X=138270 $Y=40560
X313 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=146740 51680 1 0 $X=146550 $Y=48720
X314 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=151800 40800 0 0 $X=151610 $Y=40560
X315 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=157320 73440 0 0 $X=157130 $Y=73200
X316 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=162840 73440 0 0 $X=162650 $Y=73200
X317 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=163300 57120 1 0 $X=163110 $Y=54160
X318 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=168820 57120 1 0 $X=168630 $Y=54160
X319 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=179400 35360 0 0 $X=179210 $Y=35120
X320 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=180780 68000 1 0 $X=180590 $Y=65040
X321 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=183080 40800 0 0 $X=182890 $Y=40560
X322 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=192280 51680 0 0 $X=192090 $Y=51440
X323 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=193660 57120 1 0 $X=193470 $Y=54160
X324 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=209300 51680 1 0 $X=209110 $Y=48720
X325 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=215280 73440 0 0 $X=215090 $Y=73200
X326 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=216200 62560 0 0 $X=216010 $Y=62320
X327 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=218500 51680 0 0 $X=218310 $Y=51440
X328 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=222180 57120 1 0 $X=221990 $Y=54160
X329 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=223560 40800 1 0 $X=223370 $Y=37840
X330 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=226320 62560 1 0 $X=226130 $Y=59600
X331 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=231840 62560 1 0 $X=231650 $Y=59600
X332 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=231840 73440 1 0 $X=231650 $Y=70480
X333 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235520 40800 0 0 $X=235330 $Y=40560
X334 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235520 68000 1 0 $X=235330 $Y=65040
X335 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=235980 62560 0 0 $X=235790 $Y=62320
X336 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=236440 51680 1 0 $X=236250 $Y=48720
X337 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237360 62560 1 0 $X=237170 $Y=59600
X338 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=237360 73440 1 0 $X=237170 $Y=70480
X339 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=256680 68000 1 0 $X=256490 $Y=65040
X340 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=259440 57120 1 0 $X=259250 $Y=54160
X341 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=262660 40800 1 0 $X=262470 $Y=37840
X342 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=277840 46240 1 0 $X=277650 $Y=43280
X343 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=278300 40800 1 0 $X=278110 $Y=37840
X344 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=278760 35360 0 0 $X=278570 $Y=35120
X345 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=279680 51680 1 0 $X=279490 $Y=48720
X346 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=280140 40800 0 0 $X=279950 $Y=40560
X347 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=283360 46240 1 0 $X=283170 $Y=43280
X348 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=283820 40800 1 0 $X=283630 $Y=37840
X349 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=288880 46240 1 0 $X=288690 $Y=43280
X350 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=290260 68000 1 0 $X=290070 $Y=65040
X351 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=290260 73440 1 0 $X=290070 $Y=70480
X352 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293020 40800 1 0 $X=292830 $Y=37840
X353 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=307740 57120 1 0 $X=307550 $Y=54160
X354 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=313260 57120 1 0 $X=313070 $Y=54160
X355 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=327060 62560 0 0 $X=326870 $Y=62320
X356 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=328440 68000 0 0 $X=328250 $Y=67760
X357 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=334420 68000 1 0 $X=334230 $Y=65040
X358 1 2 ICV_2 $T=19780 62560 1 0 $X=19590 $Y=59600
X359 1 2 ICV_2 $T=19780 73440 1 0 $X=19590 $Y=70480
X360 1 2 ICV_2 $T=75900 68000 1 0 $X=75710 $Y=65040
X361 1 2 ICV_2 $T=103960 40800 1 0 $X=103770 $Y=37840
X362 1 2 ICV_2 $T=103960 68000 1 0 $X=103770 $Y=65040
X363 1 2 ICV_2 $T=145820 40800 0 0 $X=145630 $Y=40560
X364 1 2 ICV_2 $T=160080 40800 1 0 $X=159890 $Y=37840
X365 1 2 ICV_2 $T=160080 78880 1 0 $X=159890 $Y=75920
X366 1 2 ICV_2 $T=188140 46240 1 0 $X=187950 $Y=43280
X367 1 2 ICV_2 $T=216200 57120 1 0 $X=216010 $Y=54160
X368 1 2 ICV_2 $T=216200 62560 1 0 $X=216010 $Y=59600
X369 1 2 ICV_2 $T=216200 78880 1 0 $X=216010 $Y=75920
X370 1 2 ICV_2 $T=230000 62560 0 0 $X=229810 $Y=62320
X371 1 2 ICV_2 $T=258060 35360 0 0 $X=257870 $Y=35120
X372 1 2 ICV_2 $T=258060 57120 0 0 $X=257870 $Y=56880
X373 1 2 ICV_2 $T=258060 62560 0 0 $X=257870 $Y=62320
X374 1 2 ICV_2 $T=258060 68000 0 0 $X=257870 $Y=67760
X375 1 2 ICV_2 $T=272320 40800 1 0 $X=272130 $Y=37840
X376 1 2 ICV_2 $T=272320 68000 1 0 $X=272130 $Y=65040
X377 1 2 ICV_2 $T=286120 40800 0 0 $X=285930 $Y=40560
X378 1 2 ICV_2 $T=286120 46240 0 0 $X=285930 $Y=46000
X379 1 2 ICV_2 $T=314180 51680 0 0 $X=313990 $Y=51440
X380 1 2 ICV_2 $T=314180 57120 0 0 $X=313990 $Y=56880
X381 1 2 ICV_2 $T=328440 57120 1 0 $X=328250 $Y=54160
X382 1 2 ICV_2 $T=328440 62560 1 0 $X=328250 $Y=59600
X383 1 2 ICV_2 $T=328440 68000 1 0 $X=328250 $Y=65040
X384 1 2 ICV_2 $T=328440 73440 1 0 $X=328250 $Y=70480
X385 1 2 ICV_2 $T=328440 78880 1 0 $X=328250 $Y=75920
X386 1 2 ICV_2 $T=342240 35360 0 0 $X=342050 $Y=35120
X387 1 2 ICV_2 $T=342240 40800 0 0 $X=342050 $Y=40560
X388 1 2 ICV_2 $T=342240 51680 0 0 $X=342050 $Y=51440
X389 1 2 ICV_2 $T=342240 57120 0 0 $X=342050 $Y=56880
X390 1 2 ICV_2 $T=342240 62560 0 0 $X=342050 $Y=62320
X391 1 2 ICV_2 $T=342240 68000 0 0 $X=342050 $Y=67760
X392 1 2 ICV_2 $T=342240 73440 0 0 $X=342050 $Y=73200
X393 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 57120 1 0 $X=17750 $Y=54160
X394 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=18400 73440 0 0 $X=18210 $Y=73200
X395 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=20240 68000 1 0 $X=20050 $Y=65040
X396 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=23920 40800 0 0 $X=23730 $Y=40560
X397 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 40800 1 0 $X=31550 $Y=37840
X398 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 51680 1 0 $X=31550 $Y=48720
X399 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=45540 46240 1 0 $X=45350 $Y=43280
X400 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 51680 1 0 $X=45810 $Y=48720
X401 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 57120 1 0 $X=45810 $Y=54160
X402 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 35360 0 0 $X=61910 $Y=35120
X403 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 57120 0 0 $X=61910 $Y=56880
X404 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=68540 78880 1 0 $X=68350 $Y=75920
X405 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73600 40800 1 0 $X=73410 $Y=37840
X406 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=90160 51680 0 0 $X=89970 $Y=51440
X407 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=101660 62560 1 0 $X=101470 $Y=59600
X408 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 40800 1 0 $X=101930 $Y=37840
X409 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 73440 1 0 $X=104230 $Y=70480
X410 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=125580 40800 0 0 $X=125390 $Y=40560
X411 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=131560 57120 0 0 $X=131370 $Y=56880
X412 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=132480 51680 1 0 $X=132290 $Y=48720
X413 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=140300 46240 0 0 $X=140110 $Y=46000
X414 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143980 40800 0 0 $X=143790 $Y=40560
X415 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=144900 78880 1 0 $X=144710 $Y=75920
X416 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=146280 62560 0 0 $X=146090 $Y=62320
X417 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=161920 46240 0 0 $X=161730 $Y=46000
X418 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=168360 51680 0 0 $X=168170 $Y=51440
X419 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=168360 73440 0 0 $X=168170 $Y=73200
X420 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174340 57120 0 0 $X=174150 $Y=56880
X421 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174340 68000 0 0 $X=174150 $Y=67760
X422 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188600 78880 1 0 $X=188410 $Y=75920
X423 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=211140 68000 0 0 $X=210950 $Y=67760
X424 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=213900 62560 1 0 $X=213710 $Y=59600
X425 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216200 40800 0 0 $X=216010 $Y=40560
X426 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 51680 1 0 $X=216470 $Y=48720
X427 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=224020 51680 0 0 $X=223830 $Y=51440
X428 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=227700 57120 1 0 $X=227510 $Y=54160
X429 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=229080 40800 1 0 $X=228890 $Y=37840
X430 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=241960 51680 1 0 $X=241770 $Y=48720
X431 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244720 73440 1 0 $X=244530 $Y=70480
X432 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=253920 73440 1 0 $X=253730 $Y=70480
X433 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 40800 0 0 $X=258330 $Y=40560
X434 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 73440 0 0 $X=258330 $Y=73200
X435 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=263580 62560 1 0 $X=263390 $Y=59600
X436 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=264040 35360 0 0 $X=263850 $Y=35120
X437 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=281980 62560 0 0 $X=281790 $Y=62320
X438 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284280 35360 0 0 $X=284090 $Y=35120
X439 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=292100 40800 0 0 $X=291910 $Y=40560
X440 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=292100 46240 0 0 $X=291910 $Y=46000
X441 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=293020 51680 1 0 $X=292830 $Y=48720
X442 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=300840 35360 0 0 $X=300650 $Y=35120
X443 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=300840 40800 1 0 $X=300650 $Y=37840
X444 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=306820 46240 0 0 $X=306630 $Y=46000
X445 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=308200 68000 0 0 $X=308010 $Y=67760
X446 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=312340 35360 0 0 $X=312150 $Y=35120
X447 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=312340 40800 0 0 $X=312150 $Y=40560
X448 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=312340 46240 0 0 $X=312150 $Y=46000
X449 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=332580 46240 1 0 $X=332390 $Y=43280
X450 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=333040 40800 0 0 $X=332850 $Y=40560
X451 1 7 sky130_fd_sc_hd__diode_2 $T=12420 46240 0 0 $X=12230 $Y=46000
X452 1 8 sky130_fd_sc_hd__diode_2 $T=39100 68000 0 0 $X=38910 $Y=67760
X453 1 369 sky130_fd_sc_hd__diode_2 $T=63940 73440 1 0 $X=63750 $Y=70480
X454 1 55 sky130_fd_sc_hd__diode_2 $T=64400 35360 0 0 $X=64210 $Y=35120
X455 1 58 sky130_fd_sc_hd__diode_2 $T=69000 73440 0 0 $X=68810 $Y=73200
X456 1 57 sky130_fd_sc_hd__diode_2 $T=70380 68000 0 0 $X=70190 $Y=67760
X457 1 372 sky130_fd_sc_hd__diode_2 $T=70840 51680 0 0 $X=70650 $Y=51440
X458 1 65 sky130_fd_sc_hd__diode_2 $T=75440 62560 0 0 $X=75250 $Y=62320
X459 1 364 sky130_fd_sc_hd__diode_2 $T=76820 46240 0 0 $X=76630 $Y=46000
X460 1 71 sky130_fd_sc_hd__diode_2 $T=79580 57120 1 0 $X=79390 $Y=54160
X461 1 8 sky130_fd_sc_hd__diode_2 $T=93840 35360 0 0 $X=93650 $Y=35120
X462 1 85 sky130_fd_sc_hd__diode_2 $T=97980 40800 0 0 $X=97790 $Y=40560
X463 1 86 sky130_fd_sc_hd__diode_2 $T=114080 73440 1 0 $X=113890 $Y=70480
X464 1 408 sky130_fd_sc_hd__diode_2 $T=120980 62560 0 0 $X=120790 $Y=62320
X465 1 87 sky130_fd_sc_hd__diode_2 $T=123280 62560 1 0 $X=123090 $Y=59600
X466 1 78 sky130_fd_sc_hd__diode_2 $T=123280 73440 0 0 $X=123090 $Y=73200
X467 1 106 sky130_fd_sc_hd__diode_2 $T=124660 73440 1 0 $X=124470 $Y=70480
X468 1 105 sky130_fd_sc_hd__diode_2 $T=125120 62560 0 0 $X=124930 $Y=62320
X469 1 106 sky130_fd_sc_hd__diode_2 $T=125120 78880 1 0 $X=124930 $Y=75920
X470 1 419 sky130_fd_sc_hd__diode_2 $T=133860 57120 0 0 $X=133670 $Y=56880
X471 1 115 sky130_fd_sc_hd__diode_2 $T=135700 62560 1 0 $X=135510 $Y=59600
X472 1 352 sky130_fd_sc_hd__diode_2 $T=138920 62560 0 0 $X=138730 $Y=62320
X473 1 117 sky130_fd_sc_hd__diode_2 $T=140760 73440 1 0 $X=140570 $Y=70480
X474 1 123 sky130_fd_sc_hd__diode_2 $T=147200 46240 0 0 $X=147010 $Y=46000
X475 1 120 sky130_fd_sc_hd__diode_2 $T=147200 68000 0 0 $X=147010 $Y=67760
X476 1 72 sky130_fd_sc_hd__diode_2 $T=148120 62560 1 0 $X=147930 $Y=59600
X477 1 426 sky130_fd_sc_hd__diode_2 $T=153180 73440 1 0 $X=152990 $Y=70480
X478 1 123 sky130_fd_sc_hd__diode_2 $T=156860 46240 0 0 $X=156670 $Y=46000
X479 1 123 sky130_fd_sc_hd__diode_2 $T=161460 46240 1 0 $X=161270 $Y=43280
X480 1 3 sky130_fd_sc_hd__diode_2 $T=164220 46240 0 0 $X=164030 $Y=46000
X481 1 352 sky130_fd_sc_hd__diode_2 $T=166520 62560 1 0 $X=166330 $Y=59600
X482 1 437 sky130_fd_sc_hd__diode_2 $T=168360 51680 1 0 $X=168170 $Y=48720
X483 1 104 sky130_fd_sc_hd__diode_2 $T=188600 35360 0 0 $X=188410 $Y=35120
X484 1 419 sky130_fd_sc_hd__diode_2 $T=191820 73440 1 0 $X=191630 $Y=70480
X485 1 157 sky130_fd_sc_hd__diode_2 $T=193200 68000 0 0 $X=193010 $Y=67760
X486 1 158 sky130_fd_sc_hd__diode_2 $T=199180 40800 1 0 $X=198990 $Y=37840
X487 1 156 sky130_fd_sc_hd__diode_2 $T=201020 51680 1 0 $X=200830 $Y=48720
X488 1 8 sky130_fd_sc_hd__diode_2 $T=208380 57120 0 0 $X=208190 $Y=56880
X489 1 459 sky130_fd_sc_hd__diode_2 $T=212520 51680 0 0 $X=212330 $Y=51440
X490 1 8 sky130_fd_sc_hd__diode_2 $T=213440 68000 0 0 $X=213250 $Y=67760
X491 1 463 sky130_fd_sc_hd__diode_2 $T=218960 51680 1 0 $X=218770 $Y=48720
X492 1 177 sky130_fd_sc_hd__diode_2 $T=221260 73440 0 0 $X=221070 $Y=73200
X493 1 451 sky130_fd_sc_hd__diode_2 $T=223100 68000 1 0 $X=222910 $Y=65040
X494 1 465 sky130_fd_sc_hd__diode_2 $T=224480 73440 1 0 $X=224290 $Y=70480
X495 1 469 sky130_fd_sc_hd__diode_2 $T=230000 57120 1 0 $X=229810 $Y=54160
X496 1 137 sky130_fd_sc_hd__diode_2 $T=237360 68000 0 0 $X=237170 $Y=67760
X497 1 193 sky130_fd_sc_hd__diode_2 $T=249320 73440 0 0 $X=249130 $Y=73200
X498 1 483 sky130_fd_sc_hd__diode_2 $T=259440 46240 0 0 $X=259250 $Y=46000
X499 1 206 sky130_fd_sc_hd__diode_2 $T=260820 73440 0 0 $X=260630 $Y=73200
X500 1 207 sky130_fd_sc_hd__diode_2 $T=261280 51680 0 0 $X=261090 $Y=51440
X501 1 487 sky130_fd_sc_hd__diode_2 $T=264040 57120 0 0 $X=263850 $Y=56880
X502 1 8 sky130_fd_sc_hd__diode_2 $T=266340 35360 0 0 $X=266150 $Y=35120
X503 1 215 sky130_fd_sc_hd__diode_2 $T=273700 78880 1 0 $X=273510 $Y=75920
X504 1 8 sky130_fd_sc_hd__diode_2 $T=294400 46240 0 0 $X=294210 $Y=46000
X505 1 228 sky130_fd_sc_hd__diode_2 $T=295780 73440 0 0 $X=295590 $Y=73200
X506 1 503 sky130_fd_sc_hd__diode_2 $T=301300 40800 0 0 $X=301110 $Y=40560
X507 1 188 sky130_fd_sc_hd__diode_2 $T=305440 62560 1 0 $X=305250 $Y=59600
X508 1 498 sky130_fd_sc_hd__diode_2 $T=305900 73440 1 0 $X=305710 $Y=70480
X509 1 231 sky130_fd_sc_hd__diode_2 $T=308660 78880 1 0 $X=308470 $Y=75920
X510 1 520 sky130_fd_sc_hd__diode_2 $T=309120 46240 0 0 $X=308930 $Y=46000
X511 1 521 sky130_fd_sc_hd__diode_2 $T=315560 40800 0 0 $X=315370 $Y=40560
X512 1 521 sky130_fd_sc_hd__diode_2 $T=315560 46240 0 0 $X=315370 $Y=46000
X513 1 459 sky130_fd_sc_hd__diode_2 $T=333040 51680 1 0 $X=332850 $Y=48720
X514 1 2 366 ICV_4 $T=58420 62560 1 0 $X=58230 $Y=59600
X515 1 2 48 ICV_4 $T=58420 62560 0 0 $X=58230 $Y=62320
X516 1 2 47 ICV_4 $T=64400 78880 1 0 $X=64210 $Y=75920
X517 1 2 61 ICV_4 $T=69460 68000 1 0 $X=69270 $Y=65040
X518 1 2 69 ICV_4 $T=77280 68000 0 0 $X=77090 $Y=67760
X519 1 2 378 ICV_4 $T=78660 57120 0 0 $X=78470 $Y=56880
X520 1 2 77 ICV_4 $T=95220 62560 0 0 $X=95030 $Y=62320
X521 1 2 356 ICV_4 $T=100280 62560 0 0 $X=100090 $Y=62320
X522 1 2 92 ICV_4 $T=109940 73440 0 0 $X=109750 $Y=73200
X523 1 2 402 ICV_4 $T=112700 51680 1 0 $X=112510 $Y=48720
X524 1 2 383 ICV_4 $T=114540 35360 0 0 $X=114350 $Y=35120
X525 1 2 407 ICV_4 $T=120520 51680 1 0 $X=120330 $Y=48720
X526 1 2 108 ICV_4 $T=128800 73440 1 0 $X=128610 $Y=70480
X527 1 2 98 ICV_4 $T=132480 73440 0 0 $X=132290 $Y=73200
X528 1 2 109 ICV_4 $T=135700 62560 0 0 $X=135510 $Y=62320
X529 1 2 388 ICV_4 $T=136160 68000 0 0 $X=135970 $Y=67760
X530 1 2 99 ICV_4 $T=137540 73440 0 0 $X=137350 $Y=73200
X531 1 2 405 ICV_4 $T=139380 51680 1 0 $X=139190 $Y=48720
X532 1 2 122 ICV_4 $T=142600 46240 0 0 $X=142410 $Y=46000
X533 1 2 120 ICV_4 $T=142600 68000 0 0 $X=142410 $Y=67760
X534 1 2 378 ICV_4 $T=144900 62560 1 0 $X=144710 $Y=59600
X535 1 2 122 ICV_4 $T=155020 57120 0 0 $X=154830 $Y=56880
X536 1 2 128 ICV_4 $T=156400 68000 0 0 $X=156210 $Y=67760
X537 1 2 329 ICV_4 $T=160540 40800 0 0 $X=160350 $Y=40560
X538 1 2 99 ICV_4 $T=161460 68000 1 0 $X=161270 $Y=65040
X539 1 2 134 ICV_4 $T=161920 57120 0 0 $X=161730 $Y=56880
X540 1 2 7 ICV_4 $T=166060 62560 0 0 $X=165870 $Y=62320
X541 1 2 410 ICV_4 $T=171580 46240 1 0 $X=171390 $Y=43280
X542 1 2 412 ICV_4 $T=176180 57120 0 0 $X=175990 $Y=56880
X543 1 2 410 ICV_4 $T=176640 51680 1 0 $X=176450 $Y=48720
X544 1 2 328 ICV_4 $T=184920 57120 1 0 $X=184730 $Y=54160
X545 1 2 438 ICV_4 $T=190440 68000 0 0 $X=190250 $Y=67760
X546 1 2 89 ICV_4 $T=193660 68000 1 0 $X=193470 $Y=65040
X547 1 2 159 ICV_4 $T=195960 73440 1 0 $X=195770 $Y=70480
X548 1 2 117 ICV_4 $T=199180 68000 1 0 $X=198990 $Y=65040
X549 1 2 162 ICV_4 $T=199640 78880 1 0 $X=199450 $Y=75920
X550 1 2 5 ICV_4 $T=202400 68000 1 0 $X=202210 $Y=65040
X551 1 2 7 ICV_4 $T=208380 73440 0 0 $X=208190 $Y=73200
X552 1 2 466 ICV_4 $T=226780 68000 0 0 $X=226590 $Y=67760
X553 1 2 475 ICV_4 $T=241040 46240 1 0 $X=240850 $Y=43280
X554 1 2 479 ICV_4 $T=247940 68000 1 0 $X=247750 $Y=65040
X555 1 2 192 ICV_4 $T=249320 57120 0 0 $X=249130 $Y=56880
X556 1 2 208 ICV_4 $T=267260 51680 0 0 $X=267070 $Y=51440
X557 1 2 169 ICV_4 $T=272320 73440 0 0 $X=272130 $Y=73200
X558 1 2 449 ICV_4 $T=273700 57120 1 0 $X=273510 $Y=54160
X559 1 2 226 ICV_4 $T=301760 46240 1 0 $X=301570 $Y=43280
X560 1 2 210 ICV_4 $T=301760 73440 0 0 $X=301570 $Y=73200
X561 1 2 236 ICV_4 $T=312340 68000 1 0 $X=312150 $Y=65040
X562 1 2 521 ICV_4 $T=319240 46240 1 0 $X=319050 $Y=43280
X563 1 2 521 ICV_4 $T=321080 40800 0 0 $X=320890 $Y=40560
X564 1 2 521 ICV_4 $T=327520 40800 0 0 $X=327330 $Y=40560
X565 1 2 525 ICV_4 $T=327520 51680 0 0 $X=327330 $Y=51440
X566 1 2 525 ICV_4 $T=330280 51680 1 0 $X=330090 $Y=48720
X567 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=27140 51680 0 0 $X=26950 $Y=51440
X568 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=31740 78880 1 0 $X=31550 $Y=75920
X569 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=36800 40800 1 0 $X=36610 $Y=37840
X570 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45540 40800 0 0 $X=45350 $Y=40560
X571 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=55660 68000 1 0 $X=55470 $Y=65040
X572 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=57960 51680 1 0 $X=57770 $Y=48720
X573 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=59800 46240 1 0 $X=59610 $Y=43280
X574 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=118220 62560 0 0 $X=118030 $Y=62320
X575 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=124200 46240 1 0 $X=124010 $Y=43280
X576 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=155020 57120 1 0 $X=154830 $Y=54160
X577 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157320 40800 0 0 $X=157130 $Y=40560
X578 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=165600 51680 1 0 $X=165410 $Y=48720
X579 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 62560 1 0 $X=185190 $Y=59600
X580 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=191360 46240 0 0 $X=191170 $Y=46000
X581 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=199180 57120 1 0 $X=198990 $Y=54160
X582 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 40800 1 0 $X=216470 $Y=37840
X583 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=220340 68000 1 0 $X=220150 $Y=65040
X584 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=221720 62560 0 0 $X=221530 $Y=62320
X585 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=240580 51680 0 0 $X=240390 $Y=51440
X586 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241040 68000 1 0 $X=240850 $Y=65040
X587 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=241500 62560 0 0 $X=241310 $Y=62320
X588 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 68000 1 0 $X=244530 $Y=65040
X589 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=253460 78880 1 0 $X=253270 $Y=75920
X590 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=255300 35360 0 0 $X=255110 $Y=35120
X591 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=258520 51680 0 0 $X=258330 $Y=51440
X592 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=262200 68000 1 0 $X=262010 $Y=65040
X593 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=271860 57120 0 0 $X=271670 $Y=56880
X594 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=278300 68000 1 0 $X=278110 $Y=65040
X595 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=287500 78880 1 0 $X=287310 $Y=75920
X596 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=295320 78880 1 0 $X=295130 $Y=75920
X597 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=295780 68000 1 0 $X=295590 $Y=65040
X598 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297160 46240 1 0 $X=296970 $Y=43280
X599 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=310960 51680 0 0 $X=310770 $Y=51440
X600 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=318780 57120 1 0 $X=318590 $Y=54160
X601 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325220 62560 1 0 $X=325030 $Y=59600
X602 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=331200 40800 1 0 $X=331010 $Y=37840
X603 1 2 34 ICV_5 $T=34960 68000 0 0 $X=34770 $Y=67760
X604 1 2 75 ICV_5 $T=81880 73440 0 0 $X=81690 $Y=73200
X605 1 2 395 ICV_5 $T=105340 62560 0 0 $X=105150 $Y=62320
X606 1 2 88 ICV_5 $T=105340 78880 1 0 $X=105150 $Y=75920
X607 1 2 98 ICV_5 $T=120980 73440 1 0 $X=120790 $Y=70480
X608 1 2 416 ICV_5 $T=137080 68000 1 0 $X=136890 $Y=65040
X609 1 2 405 ICV_5 $T=138460 46240 1 0 $X=138270 $Y=43280
X610 1 2 415 ICV_5 $T=139840 51680 0 0 $X=139650 $Y=51440
X611 1 2 425 ICV_5 $T=157780 51680 0 0 $X=157590 $Y=51440
X612 1 2 445 ICV_5 $T=174340 57120 1 0 $X=174150 $Y=54160
X613 1 2 128 ICV_5 $T=233680 68000 0 0 $X=233490 $Y=67760
X614 1 2 186 ICV_5 $T=240120 78880 1 0 $X=239930 $Y=75920
X615 1 2 187 ICV_5 $T=245180 73440 0 0 $X=244990 $Y=73200
X616 1 2 191 ICV_5 $T=247020 73440 1 0 $X=246830 $Y=70480
X617 1 2 8 ICV_5 $T=252540 46240 0 0 $X=252350 $Y=46000
X618 1 2 489 ICV_5 $T=265880 57120 1 0 $X=265690 $Y=54160
X619 1 2 491 ICV_5 $T=268640 40800 1 0 $X=268450 $Y=37840
X620 1 2 512 ICV_5 $T=301760 62560 1 0 $X=301570 $Y=59600
X621 1 2 246 ICV_5 $T=338100 35360 0 0 $X=337910 $Y=35120
X622 1 2 248 ICV_5 $T=338100 68000 0 0 $X=337910 $Y=67760
X623 1 2 249 ICV_5 $T=338560 40800 0 0 $X=338370 $Y=40560
X624 1 2 250 ICV_5 $T=338560 57120 0 0 $X=338370 $Y=56880
X625 1 2 245 ICV_5 $T=338560 73440 0 0 $X=338370 $Y=73200
X626 1 2 9 ICV_6 $T=7820 46240 0 0 $X=7630 $Y=46000
X627 1 2 8 ICV_6 $T=14260 46240 1 0 $X=14070 $Y=43280
X628 1 2 15 ICV_6 $T=14260 51680 1 0 $X=14070 $Y=48720
X629 1 2 23 ICV_6 $T=23920 35360 0 0 $X=23730 $Y=35120
X630 1 2 350 ICV_6 $T=34040 68000 1 0 $X=33850 $Y=65040
X631 1 2 37 ICV_6 $T=46460 35360 0 0 $X=46270 $Y=35120
X632 1 2 360 ICV_6 $T=51520 57120 1 0 $X=51330 $Y=54160
X633 1 2 47 ICV_6 $T=55200 78880 1 0 $X=55010 $Y=75920
X634 1 2 46 ICV_6 $T=55660 35360 0 0 $X=55470 $Y=35120
X635 1 2 389 ICV_6 $T=98440 51680 1 0 $X=98250 $Y=48720
X636 1 2 90 ICV_6 $T=109020 73440 1 0 $X=108830 $Y=70480
X637 1 2 399 ICV_6 $T=110400 57120 0 0 $X=110210 $Y=56880
X638 1 2 78 ICV_6 $T=120060 78880 1 0 $X=119870 $Y=75920
X639 1 2 413 ICV_6 $T=127420 51680 1 0 $X=127230 $Y=48720
X640 1 2 132 ICV_6 $T=163300 40800 0 0 $X=163110 $Y=40560
X641 1 2 137 ICV_6 $T=168360 68000 1 0 $X=168170 $Y=65040
X642 1 2 123 ICV_6 $T=169280 35360 0 0 $X=169090 $Y=35120
X643 1 2 148 ICV_6 $T=184000 51680 0 0 $X=183810 $Y=51440
X644 1 2 457 ICV_6 $T=210680 46240 1 0 $X=210490 $Y=43280
X645 1 2 472 ICV_6 $T=235520 46240 1 0 $X=235330 $Y=43280
X646 1 2 480 ICV_6 $T=248400 46240 1 0 $X=248210 $Y=43280
X647 1 2 196 ICV_6 $T=276920 68000 0 0 $X=276730 $Y=67760
X648 1 2 493 ICV_6 $T=281060 46240 0 0 $X=280870 $Y=46000
X649 1 2 498 ICV_6 $T=293020 62560 1 0 $X=292830 $Y=59600
X650 1 2 504 ICV_6 $T=296240 40800 0 0 $X=296050 $Y=40560
X651 1 2 511 ICV_6 $T=302680 57120 0 0 $X=302490 $Y=56880
X652 1 2 504 ICV_6 $T=316940 40800 1 0 $X=316750 $Y=37840
X653 1 2 524 ICV_6 $T=323380 73440 1 0 $X=323190 $Y=70480
X654 1 2 8 ICV_6 $T=343620 46240 0 0 $X=343430 $Y=46000
X655 1 7 8 ICV_7 $T=7820 40800 1 0 $X=7630 $Y=37840
X656 1 7 8 ICV_7 $T=7820 57120 1 0 $X=7630 $Y=54160
X657 1 7 12 ICV_7 $T=7820 62560 1 0 $X=7630 $Y=59600
X658 1 7 8 ICV_7 $T=7820 73440 1 0 $X=7630 $Y=70480
X659 1 7 14 ICV_7 $T=7820 78880 1 0 $X=7630 $Y=75920
X660 1 343 8 ICV_7 $T=15640 68000 0 0 $X=15450 $Y=67760
X661 1 7 8 ICV_7 $T=20240 35360 0 0 $X=20050 $Y=35120
X662 1 8 22 ICV_7 $T=20240 73440 0 0 $X=20050 $Y=73200
X663 1 8 344 ICV_7 $T=22540 62560 0 0 $X=22350 $Y=62320
X664 1 8 345 ICV_7 $T=24380 51680 0 0 $X=24190 $Y=51440
X665 1 26 7 ICV_7 $T=25760 40800 0 0 $X=25570 $Y=40560
X666 1 27 347 ICV_7 $T=28060 46240 0 0 $X=27870 $Y=46000
X667 1 346 349 ICV_7 $T=28060 57120 0 0 $X=27870 $Y=56880
X668 1 8 351 ICV_7 $T=34040 40800 1 0 $X=33850 $Y=37840
X669 1 39 356 ICV_7 $T=43700 51680 0 0 $X=43510 $Y=51440
X670 1 353 39 ICV_7 $T=44160 57120 0 0 $X=43970 $Y=56880
X671 1 42 39 ICV_7 $T=46460 62560 0 0 $X=46270 $Y=62320
X672 1 356 43 ICV_7 $T=47840 73440 0 0 $X=47650 $Y=73200
X673 1 8 359 ICV_7 $T=48300 40800 0 0 $X=48110 $Y=40560
X674 1 358 329 ICV_7 $T=49220 62560 1 0 $X=49030 $Y=59600
X675 1 39 42 ICV_7 $T=51520 78880 1 0 $X=51330 $Y=75920
X676 1 7 8 ICV_7 $T=51980 35360 0 0 $X=51790 $Y=35120
X677 1 39 42 ICV_7 $T=52440 68000 0 0 $X=52250 $Y=67760
X678 1 362 36 ICV_7 $T=54740 62560 0 0 $X=54550 $Y=62320
X679 1 363 48 ICV_7 $T=55200 51680 0 0 $X=55010 $Y=51440
X680 1 45 365 ICV_7 $T=56120 68000 0 0 $X=55930 $Y=67760
X681 1 368 45 ICV_7 $T=60260 73440 1 0 $X=60070 $Y=70480
X682 1 51 54 ICV_7 $T=60720 78880 1 0 $X=60530 $Y=75920
X683 1 51 371 ICV_7 $T=63020 51680 1 0 $X=62830 $Y=48720
X684 1 353 57 ICV_7 $T=64400 57120 1 0 $X=64210 $Y=54160
X685 1 49 49 ICV_7 $T=65320 73440 0 0 $X=65130 $Y=73200
X686 1 58 57 ICV_7 $T=65780 68000 1 0 $X=65590 $Y=65040
X687 1 48 372 ICV_7 $T=68080 57120 1 0 $X=67890 $Y=54160
X688 1 373 375 ICV_7 $T=69460 46240 0 0 $X=69270 $Y=46000
X689 1 65 56 ICV_7 $T=72220 68000 1 0 $X=72030 $Y=65040
X690 1 377 377 ICV_7 $T=73140 46240 0 0 $X=72950 $Y=46000
X691 1 375 381 ICV_7 $T=77280 40800 1 0 $X=77090 $Y=37840
X692 1 69 56 ICV_7 $T=78200 73440 0 0 $X=78010 $Y=73200
X693 1 70 381 ICV_7 $T=79120 35360 0 0 $X=78930 $Y=35120
X694 1 61 385 ICV_7 $T=82340 62560 1 0 $X=82150 $Y=59600
X695 1 386 69 ICV_7 $T=85560 73440 0 0 $X=85370 $Y=73200
X696 1 387 389 ICV_7 $T=86020 62560 1 0 $X=85830 $Y=59600
X697 1 385 71 ICV_7 $T=89700 51680 1 0 $X=89510 $Y=48720
X698 1 65 77 ICV_7 $T=91540 68000 0 0 $X=91350 $Y=67760
X699 1 375 391 ICV_7 $T=92000 46240 1 0 $X=91810 $Y=43280
X700 1 70 81 ICV_7 $T=95220 46240 0 0 $X=95030 $Y=46000
X701 1 377 67 ICV_7 $T=95220 57120 0 0 $X=95030 $Y=56880
X702 1 78 389 ICV_7 $T=95220 68000 1 0 $X=95030 $Y=65040
X703 1 393 8 ICV_7 $T=99820 51680 0 0 $X=99630 $Y=51440
X704 1 86 87 ICV_7 $T=101200 73440 0 0 $X=101010 $Y=73200
X705 1 383 374 ICV_7 $T=103500 46240 0 0 $X=103310 $Y=46000
X706 1 49 383 ICV_7 $T=106720 57120 0 0 $X=106530 $Y=56880
X707 1 398 69 ICV_7 $T=109020 62560 0 0 $X=108830 $Y=62320
X708 1 400 381 ICV_7 $T=110860 35360 0 0 $X=110670 $Y=35120
X709 1 401 403 ICV_7 $T=111320 40800 0 0 $X=111130 $Y=40560
X710 1 94 92 ICV_7 $T=111780 46240 0 0 $X=111590 $Y=46000
X711 1 405 409 ICV_7 $T=121440 68000 0 0 $X=121250 $Y=67760
X712 1 92 411 ICV_7 $T=123280 46240 0 0 $X=123090 $Y=46000
X713 1 410 412 ICV_7 $T=123740 57120 0 0 $X=123550 $Y=56880
X714 1 405 398 ICV_7 $T=125120 68000 0 0 $X=124930 $Y=67760
X715 1 110 111 ICV_7 $T=127880 40800 0 0 $X=127690 $Y=40560
X716 1 405 412 ICV_7 $T=131100 51680 0 0 $X=130910 $Y=51440
X717 1 414 113 ICV_7 $T=133400 57120 1 0 $X=133210 $Y=54160
X718 1 105 114 ICV_7 $T=133400 68000 1 0 $X=133210 $Y=65040
X719 1 419 115 ICV_7 $T=137540 57120 1 0 $X=137350 $Y=54160
X720 1 101 422 ICV_7 $T=138460 35360 0 0 $X=138270 $Y=35120
X721 1 87 113 ICV_7 $T=138920 68000 0 0 $X=138730 $Y=67760
X722 1 423 424 ICV_7 $T=141220 68000 1 0 $X=141030 $Y=65040
X723 1 118 127 ICV_7 $T=147200 73440 0 0 $X=147010 $Y=73200
X724 1 124 116 ICV_7 $T=147200 78880 1 0 $X=147010 $Y=75920
X725 1 414 128 ICV_7 $T=148120 57120 1 0 $X=147930 $Y=54160
X726 1 72 129 ICV_7 $T=148120 62560 0 0 $X=147930 $Y=62320
X727 1 427 99 ICV_7 $T=149500 73440 1 0 $X=149310 $Y=70480
X728 1 3 433 ICV_7 $T=153180 46240 0 0 $X=152990 $Y=46000
X729 1 429 428 ICV_7 $T=154100 51680 0 0 $X=153910 $Y=51440
X730 1 138 140 ICV_7 $T=166060 78880 1 0 $X=165870 $Y=75920
X731 1 132 437 ICV_7 $T=168360 40800 0 0 $X=168170 $Y=40560
X732 1 112 127 ICV_7 $T=169740 78880 1 0 $X=169550 $Y=75920
X733 1 441 443 ICV_7 $T=171580 40800 1 0 $X=171390 $Y=37840
X734 1 435 444 ICV_7 $T=172040 73440 1 0 $X=171850 $Y=70480
X735 1 395 129 ICV_7 $T=174340 68000 1 0 $X=174150 $Y=65040
X736 1 144 378 ICV_7 $T=175260 40800 1 0 $X=175070 $Y=37840
X737 1 434 149 ICV_7 $T=178020 68000 1 0 $X=177830 $Y=65040
X738 1 330 3 ICV_7 $T=178940 57120 0 0 $X=178750 $Y=56880
X739 1 137 434 ICV_7 $T=179400 62560 0 0 $X=179210 $Y=62320
X740 1 329 330 ICV_7 $T=180320 40800 0 0 $X=180130 $Y=40560
X741 1 145 395 ICV_7 $T=180320 51680 0 0 $X=180130 $Y=51440
X742 1 329 4 ICV_7 $T=182620 62560 1 0 $X=182430 $Y=59600
X743 1 151 152 ICV_7 $T=182620 73440 1 0 $X=182430 $Y=70480
X744 1 427 150 ICV_7 $T=184000 73440 0 0 $X=183810 $Y=73200
X745 1 153 154 ICV_7 $T=184920 35360 0 0 $X=184730 $Y=35120
X746 1 149 419 ICV_7 $T=188140 62560 0 0 $X=187950 $Y=62320
X747 1 8 447 ICV_7 $T=188600 46240 0 0 $X=188410 $Y=46000
X748 1 6 334 ICV_7 $T=189520 51680 0 0 $X=189330 $Y=51440
X749 1 452 454 ICV_7 $T=194580 46240 0 0 $X=194390 $Y=46000
X750 1 158 154 ICV_7 $T=195500 40800 0 0 $X=195310 $Y=40560
X751 1 331 456 ICV_7 $T=203780 62560 1 0 $X=203590 $Y=59600
X752 1 5 4 ICV_7 $T=209760 68000 1 0 $X=209570 $Y=65040
X753 1 461 173 ICV_7 $T=217120 35360 0 0 $X=216930 $Y=35120
X754 1 460 464 ICV_7 $T=217580 68000 1 0 $X=217390 $Y=65040
X755 1 462 175 ICV_7 $T=218500 40800 0 0 $X=218310 $Y=40560
X756 1 178 463 ICV_7 $T=222180 40800 0 0 $X=221990 $Y=40560
X757 1 139 180 ICV_7 $T=222180 46240 0 0 $X=221990 $Y=46000
X758 1 178 175 ICV_7 $T=228160 46240 1 0 $X=227970 $Y=43280
X759 1 173 473 ICV_7 $T=231380 35360 0 0 $X=231190 $Y=35120
X760 1 471 178 ICV_7 $T=231840 46240 1 0 $X=231650 $Y=43280
X761 1 180 180 ICV_7 $T=237820 51680 0 0 $X=237630 $Y=51440
X762 1 474 466 ICV_7 $T=239200 57120 0 0 $X=239010 $Y=56880
X763 1 474 115 ICV_7 $T=243800 51680 0 0 $X=243610 $Y=51440
X764 1 466 477 ICV_7 $T=244260 62560 0 0 $X=244070 $Y=62320
X765 1 197 199 ICV_7 $T=250700 78880 1 0 $X=250510 $Y=75920
X766 1 8 192 ICV_7 $T=254380 57120 0 0 $X=254190 $Y=56880
X767 1 137 456 ICV_7 $T=254380 62560 0 0 $X=254190 $Y=62320
X768 1 484 195 ICV_7 $T=259900 40800 1 0 $X=259710 $Y=37840
X769 1 169 486 ICV_7 $T=263120 73440 1 0 $X=262930 $Y=70480
X770 1 481 487 ICV_7 $T=264960 46240 1 0 $X=264770 $Y=43280
X771 1 210 211 ICV_7 $T=264960 62560 0 0 $X=264770 $Y=62320
X772 1 157 213 ICV_7 $T=268180 78880 1 0 $X=267990 $Y=75920
X773 1 53 495 ICV_7 $T=274620 57120 0 0 $X=274430 $Y=56880
X774 1 191 218 ICV_7 $T=276460 57120 1 0 $X=276270 $Y=54160
X775 1 216 216 ICV_7 $T=276920 62560 0 0 $X=276730 $Y=62320
X776 1 488 492 ICV_7 $T=277380 46240 0 0 $X=277190 $Y=46000
X777 1 8 496 ICV_7 $T=280600 51680 0 0 $X=280410 $Y=51440
X778 1 215 194 ICV_7 $T=280600 73440 0 0 $X=280410 $Y=73200
X779 1 495 177 ICV_7 $T=287500 68000 1 0 $X=287310 $Y=65040
X780 1 8 224 ICV_7 $T=290260 40800 1 0 $X=290070 $Y=37840
X781 1 223 186 ICV_7 $T=290260 78880 1 0 $X=290070 $Y=75920
X782 1 495 483 ICV_7 $T=293940 57120 0 0 $X=293750 $Y=56880
X783 1 226 506 ICV_7 $T=294860 51680 1 0 $X=294670 $Y=48720
X784 1 342 507 ICV_7 $T=294860 68000 0 0 $X=294670 $Y=67760
X785 1 177 510 ICV_7 $T=297160 62560 0 0 $X=296970 $Y=62320
X786 1 230 221 ICV_7 $T=298540 68000 0 0 $X=298350 $Y=67760
X787 1 513 514 ICV_7 $T=302220 68000 1 0 $X=302030 $Y=65040
X788 1 515 235 ICV_7 $T=304980 46240 1 0 $X=304790 $Y=43280
X789 1 498 514 ICV_7 $T=307740 62560 0 0 $X=307550 $Y=62320
X790 1 483 498 ICV_7 $T=308200 51680 0 0 $X=308010 $Y=51440
X791 1 498 522 ICV_7 $T=314640 73440 1 0 $X=314450 $Y=70480
X792 1 7 8 ICV_7 $T=334420 35360 0 0 $X=334230 $Y=35120
X793 1 7 8 ICV_7 $T=334420 51680 0 0 $X=334230 $Y=51440
X794 1 7 8 ICV_7 $T=334420 68000 0 0 $X=334230 $Y=67760
X795 1 7 8 ICV_7 $T=334880 40800 0 0 $X=334690 $Y=40560
X796 1 7 8 ICV_7 $T=334880 57120 0 0 $X=334690 $Y=56880
X797 1 7 8 ICV_7 $T=334880 73440 0 0 $X=334690 $Y=73200
X798 1 247 520 ICV_7 $T=338100 51680 0 0 $X=337910 $Y=51440
X799 1 2 7 10 8 2 16 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 40800 0 0 $X=7630 $Y=40560
X800 1 2 7 9 8 2 17 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 51680 0 0 $X=7630 $Y=51440
X801 1 2 7 11 8 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 57120 0 0 $X=7630 $Y=56880
X802 1 2 7 12 8 2 19 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 62560 0 0 $X=7630 $Y=62320
X803 1 2 7 342 8 2 20 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 73440 0 0 $X=7630 $Y=73200
X804 1 2 7 13 8 2 21 1 sky130_fd_sc_hd__dfrtp_4 $T=8280 35360 0 0 $X=8090 $Y=35120
X805 1 2 7 15 8 2 25 1 sky130_fd_sc_hd__dfrtp_4 $T=14260 46240 0 0 $X=14070 $Y=46000
X806 1 2 526 343 8 2 28 1 sky130_fd_sc_hd__dfrtp_4 $T=19320 68000 0 0 $X=19130 $Y=67760
X807 1 2 7 23 8 2 30 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 40800 1 0 $X=20970 $Y=37840
X808 1 2 7 24 8 2 31 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 51680 1 0 $X=20970 $Y=48720
X809 1 2 527 22 8 2 32 1 sky130_fd_sc_hd__dfrtp_4 $T=21160 78880 1 0 $X=20970 $Y=75920
X810 1 2 528 344 8 2 34 1 sky130_fd_sc_hd__dfrtp_4 $T=22540 68000 1 0 $X=22350 $Y=65040
X811 1 2 529 345 8 2 33 1 sky130_fd_sc_hd__dfrtp_4 $T=24380 57120 1 0 $X=24190 $Y=54160
X812 1 2 7 26 8 2 35 1 sky130_fd_sc_hd__dfrtp_4 $T=27600 46240 1 0 $X=27410 $Y=43280
X813 1 2 7 29 8 2 40 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 35360 0 0 $X=34770 $Y=35120
X814 1 2 530 351 8 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 40800 0 0 $X=34770 $Y=40560
X815 1 2 7 27 8 2 41 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 46240 0 0 $X=34770 $Y=46000
X816 1 2 531 354 8 2 43 1 sky130_fd_sc_hd__dfrtp_4 $T=40940 68000 0 0 $X=40750 $Y=67760
X817 1 2 532 359 8 2 50 1 sky130_fd_sc_hd__dfrtp_4 $T=49220 46240 1 0 $X=49030 $Y=43280
X818 1 2 7 46 8 2 52 1 sky130_fd_sc_hd__dfrtp_4 $T=51980 40800 1 0 $X=51790 $Y=37840
X819 1 2 533 392 8 2 85 1 sky130_fd_sc_hd__dfrtp_4 $T=95680 35360 0 0 $X=95490 $Y=35120
X820 1 2 534 393 8 2 96 1 sky130_fd_sc_hd__dfrtp_4 $T=103500 51680 0 0 $X=103310 $Y=51440
X821 1 2 535 103 8 2 111 1 sky130_fd_sc_hd__dfrtp_4 $T=121440 35360 0 0 $X=121250 $Y=35120
X822 1 2 536 135 8 2 123 1 sky130_fd_sc_hd__dfrtp_4 $T=157780 35360 0 0 $X=157590 $Y=35120
X823 1 2 537 447 8 2 3 1 sky130_fd_sc_hd__dfrtp_4 $T=189520 51680 1 0 $X=189330 $Y=48720
X824 1 2 538 338 8 2 176 1 sky130_fd_sc_hd__dfrtp_4 $T=210220 57120 0 0 $X=210030 $Y=56880
X825 1 2 539 457 8 2 459 1 sky130_fd_sc_hd__dfrtp_4 $T=210680 46240 0 0 $X=210490 $Y=46000
X826 1 2 540 460 8 2 120 1 sky130_fd_sc_hd__dfrtp_4 $T=215280 68000 0 0 $X=215090 $Y=67760
X827 1 2 541 467 8 2 130 1 sky130_fd_sc_hd__dfrtp_4 $T=224940 68000 1 0 $X=224750 $Y=65040
X828 1 2 542 185 8 2 190 1 sky130_fd_sc_hd__dfrtp_4 $T=237360 35360 0 0 $X=237170 $Y=35120
X829 1 2 543 475 8 2 192 1 sky130_fd_sc_hd__dfrtp_4 $T=241040 46240 0 0 $X=240850 $Y=46000
X830 1 2 544 480 8 2 7 1 sky130_fd_sc_hd__dfrtp_4 $T=248400 51680 1 0 $X=248210 $Y=48720
X831 1 2 545 478 8 2 196 1 sky130_fd_sc_hd__dfrtp_4 $T=253000 62560 1 0 $X=252810 $Y=59600
X832 1 2 546 212 8 2 207 1 sky130_fd_sc_hd__dfrtp_4 $T=268180 35360 0 0 $X=267990 $Y=35120
X833 1 2 547 496 8 2 218 1 sky130_fd_sc_hd__dfrtp_4 $T=280600 57120 1 0 $X=280410 $Y=54160
X834 1 2 7 224 8 2 232 1 sky130_fd_sc_hd__dfrtp_4 $T=290260 35360 0 0 $X=290070 $Y=35120
X835 1 2 548 505 8 2 226 1 sky130_fd_sc_hd__dfrtp_4 $T=296240 46240 0 0 $X=296050 $Y=46000
X836 1 2 549 519 8 2 342 1 sky130_fd_sc_hd__dfrtp_4 $T=307280 62560 1 0 $X=307090 $Y=59600
X837 1 2 550 524 8 2 245 1 sky130_fd_sc_hd__dfrtp_4 $T=323380 73440 0 0 $X=323190 $Y=73200
X838 1 2 7 246 8 2 251 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 40800 1 0 $X=334230 $Y=37840
X839 1 2 7 247 8 2 252 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 57120 1 0 $X=334230 $Y=54160
X840 1 2 7 248 8 2 253 1 sky130_fd_sc_hd__dfrtp_4 $T=334420 73440 1 0 $X=334230 $Y=70480
X841 1 2 7 249 8 2 254 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 46240 1 0 $X=334690 $Y=43280
X842 1 2 7 459 8 2 255 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 51680 1 0 $X=334690 $Y=48720
X843 1 2 7 250 8 2 256 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 62560 1 0 $X=334690 $Y=59600
X844 1 2 7 245 8 2 257 1 sky130_fd_sc_hd__dfrtp_4 $T=334880 78880 1 0 $X=334690 $Y=75920
X845 1 2 24 ICV_12 $T=25760 46240 0 0 $X=25570 $Y=46000
X846 1 2 8 ICV_12 $T=29440 40800 0 0 $X=29250 $Y=40560
X847 1 2 8 ICV_12 $T=34040 51680 1 0 $X=33850 $Y=48720
X848 1 2 53 ICV_12 $T=65320 62560 0 0 $X=65130 $Y=62320
X849 1 2 385 ICV_12 $T=87400 51680 1 0 $X=87210 $Y=48720
X850 1 2 394 ICV_12 $T=101660 57120 1 0 $X=101470 $Y=54160
X851 1 2 96 ICV_12 $T=115460 46240 0 0 $X=115270 $Y=46000
X852 1 2 399 ICV_12 $T=118220 57120 1 0 $X=118030 $Y=54160
X853 1 2 395 ICV_12 $T=121440 57120 0 0 $X=121250 $Y=56880
X854 1 2 412 ICV_12 $T=133400 62560 0 0 $X=133210 $Y=62320
X855 1 2 95 ICV_12 $T=134780 51680 1 0 $X=134590 $Y=48720
X856 1 2 434 ICV_12 $T=157780 57120 1 0 $X=157590 $Y=54160
X857 1 2 432 ICV_12 $T=157780 62560 1 0 $X=157590 $Y=59600
X858 1 2 395 ICV_12 $T=189520 62560 1 0 $X=189330 $Y=59600
X859 1 2 153 ICV_12 $T=197800 35360 0 0 $X=197610 $Y=35120
X860 1 2 449 ICV_12 $T=199180 62560 1 0 $X=198990 $Y=59600
X861 1 2 183 ICV_12 $T=230460 78880 1 0 $X=230270 $Y=75920
X862 1 2 165 ICV_12 $T=235520 73440 0 0 $X=235330 $Y=73200
X863 1 2 494 ICV_12 $T=270020 57120 1 0 $X=269830 $Y=54160
X864 1 2 202 ICV_12 $T=281980 68000 0 0 $X=281790 $Y=67760
X865 1 2 357 ICV_13 $T=44160 68000 1 0 $X=43970 $Y=65040
X866 1 2 370 ICV_13 $T=62560 62560 1 0 $X=62370 $Y=59600
X867 1 2 63 ICV_13 $T=70380 35360 0 0 $X=70190 $Y=35120
X868 1 2 57 ICV_13 $T=70840 57120 0 0 $X=70650 $Y=56880
X869 1 2 379 ICV_13 $T=72220 46240 1 0 $X=72030 $Y=43280
X870 1 2 362 ICV_13 $T=76360 51680 1 0 $X=76170 $Y=48720
X871 1 2 77 ICV_13 $T=86020 57120 0 0 $X=85830 $Y=56880
X872 1 2 64 ICV_13 $T=87400 68000 1 0 $X=87210 $Y=65040
X873 1 2 369 ICV_13 $T=87860 57120 1 0 $X=87670 $Y=54160
X874 1 2 51 ICV_13 $T=97980 57120 0 0 $X=97790 $Y=56880
X875 1 2 374 ICV_13 $T=104420 57120 1 0 $X=104230 $Y=54160
X876 1 2 92 ICV_13 $T=114080 51680 0 0 $X=113890 $Y=51440
X877 1 2 403 ICV_13 $T=121440 46240 1 0 $X=121250 $Y=43280
X878 1 2 112 ICV_13 $T=128340 78880 1 0 $X=128150 $Y=75920
X879 1 2 113 ICV_13 $T=133400 46240 0 0 $X=133210 $Y=46000
X880 1 2 126 ICV_13 $T=146280 35360 0 0 $X=146090 $Y=35120
X881 1 2 412 ICV_13 $T=146280 57120 0 0 $X=146090 $Y=56880
X882 1 2 8 ICV_13 $T=154100 35360 0 0 $X=153910 $Y=35120
X883 1 2 434 ICV_13 $T=156400 51680 1 0 $X=156210 $Y=48720
X884 1 2 120 ICV_13 $T=158240 62560 0 0 $X=158050 $Y=62320
X885 1 2 353 ICV_13 $T=172500 62560 1 0 $X=172310 $Y=59600
X886 1 2 5 ICV_13 $T=181700 68000 0 0 $X=181510 $Y=67760
X887 1 2 446 ICV_13 $T=188600 40800 0 0 $X=188410 $Y=40560
X888 1 2 159 ICV_13 $T=203320 73440 1 0 $X=203130 $Y=70480
X889 1 2 458 ICV_13 $T=212520 68000 1 0 $X=212330 $Y=65040
X890 1 2 6 ICV_13 $T=212520 73440 1 0 $X=212330 $Y=70480
X891 1 2 182 ICV_13 $T=226320 51680 1 0 $X=226130 $Y=48720
X892 1 2 470 ICV_13 $T=226320 73440 0 0 $X=226130 $Y=73200
X893 1 2 152 ICV_13 $T=234140 78880 1 0 $X=233950 $Y=75920
X894 1 2 470 ICV_13 $T=243340 68000 0 0 $X=243150 $Y=67760
X895 1 2 203 ICV_13 $T=256220 46240 1 0 $X=256030 $Y=43280
X896 1 2 485 ICV_13 $T=258980 51680 1 0 $X=258790 $Y=48720
X897 1 2 169 ICV_13 $T=259440 78880 1 0 $X=259250 $Y=75920
X898 1 2 210 ICV_13 $T=264040 68000 0 0 $X=263850 $Y=67760
X899 1 2 490 ICV_13 $T=264960 40800 0 0 $X=264770 $Y=40560
X900 1 2 187 ICV_13 $T=265880 73440 1 0 $X=265690 $Y=70480
X901 1 2 483 ICV_13 $T=267260 46240 0 0 $X=267070 $Y=46000
X902 1 2 492 ICV_13 $T=268180 51680 1 0 $X=267990 $Y=48720
X903 1 2 196 ICV_13 $T=270940 68000 0 0 $X=270750 $Y=67760
X904 1 2 194 ICV_13 $T=276920 78880 1 0 $X=276730 $Y=75920
X905 1 2 221 ICV_13 $T=282440 57120 0 0 $X=282250 $Y=56880
X906 1 2 497 ICV_13 $T=282440 62560 1 0 $X=282250 $Y=59600
X907 1 2 198 ICV_13 $T=284740 78880 1 0 $X=284550 $Y=75920
X908 1 2 7 ICV_13 $T=286580 35360 0 0 $X=286390 $Y=35120
X909 1 2 505 ICV_13 $T=294400 46240 1 0 $X=294210 $Y=43280
X910 1 2 221 ICV_13 $T=298080 51680 0 0 $X=297890 $Y=51440
X911 1 2 518 ICV_13 $T=310500 62560 0 0 $X=310310 $Y=62320
X912 1 2 241 ICV_13 $T=310500 73440 0 0 $X=310310 $Y=73200
X913 1 2 525 ICV_13 $T=318320 51680 1 0 $X=318130 $Y=48720
X914 1 2 8 ICV_13 $T=319700 73440 0 0 $X=319510 $Y=73200
X915 1 2 521 ICV_13 $T=320160 51680 0 0 $X=319970 $Y=51440
X916 1 2 525 ICV_13 $T=324760 51680 1 0 $X=324570 $Y=48720
X917 1 8 ICV_15 $T=31740 40800 0 0 $X=31550 $Y=40560
X918 1 7 ICV_15 $T=31740 46240 0 0 $X=31550 $Y=46000
X919 1 33 ICV_15 $T=31740 57120 0 0 $X=31550 $Y=56880
X920 1 349 ICV_15 $T=31740 62560 0 0 $X=31550 $Y=62320
X921 1 48 ICV_15 $T=59800 68000 0 0 $X=59610 $Y=67760
X922 1 71 ICV_15 $T=87860 62560 0 0 $X=87670 $Y=62320
X923 1 99 ICV_15 $T=115920 57120 0 0 $X=115730 $Y=56880
X924 1 425 ICV_15 $T=143980 51680 0 0 $X=143790 $Y=51440
X925 1 134 ICV_15 $T=158240 46240 1 0 $X=158050 $Y=43280
X926 1 3 ICV_15 $T=172040 40800 0 0 $X=171850 $Y=40560
X927 1 140 ICV_15 $T=186300 68000 1 0 $X=186110 $Y=65040
X928 1 118 ICV_15 $T=186300 73440 1 0 $X=186110 $Y=70480
X929 1 160 ICV_15 $T=200100 35360 0 0 $X=199910 $Y=35120
X930 1 145 ICV_15 $T=200100 73440 0 0 $X=199910 $Y=73200
X931 1 476 ICV_15 $T=242420 57120 1 0 $X=242230 $Y=54160
X932 1 482 ICV_15 $T=256220 40800 0 0 $X=256030 $Y=40560
X933 1 188 ICV_15 $T=256220 46240 0 0 $X=256030 $Y=46000
X934 1 499 ICV_15 $T=284280 51680 0 0 $X=284090 $Y=51440
X935 1 500 ICV_15 $T=284280 62560 0 0 $X=284090 $Y=62320
X936 1 222 ICV_15 $T=284280 68000 0 0 $X=284090 $Y=67760
X937 1 219 ICV_15 $T=284280 73440 0 0 $X=284090 $Y=73200
X938 1 503 ICV_15 $T=298540 40800 1 0 $X=298350 $Y=37840
X939 1 508 ICV_15 $T=298540 51680 1 0 $X=298350 $Y=48720
X940 1 510 ICV_15 $T=298540 57120 1 0 $X=298350 $Y=54160
X941 1 177 ICV_15 $T=298540 68000 1 0 $X=298350 $Y=65040
X942 1 229 ICV_15 $T=298540 78880 1 0 $X=298350 $Y=75920
X943 1 2 8 ICV_16 $T=7820 68000 1 0 $X=7630 $Y=65040
X944 1 2 342 ICV_16 $T=7820 68000 0 0 $X=7630 $Y=67760
X945 1 2 11 ICV_16 $T=11500 57120 1 0 $X=11310 $Y=54160
X946 1 2 28 ICV_16 $T=34960 73440 0 0 $X=34770 $Y=73200
X947 1 2 349 ICV_16 $T=39100 46240 1 0 $X=38910 $Y=43280
X948 1 2 354 ICV_16 $T=40940 73440 1 0 $X=40750 $Y=70480
X949 1 2 50 ICV_16 $T=63020 40800 0 0 $X=62830 $Y=40560
X950 1 2 356 ICV_16 $T=63020 46240 0 0 $X=62830 $Y=46000
X951 1 2 73 ICV_16 $T=79580 73440 1 0 $X=79390 $Y=70480
X952 1 2 378 ICV_16 $T=81420 62560 0 0 $X=81230 $Y=62320
X953 1 2 72 ICV_16 $T=82340 68000 0 0 $X=82150 $Y=67760
X954 1 2 388 ICV_16 $T=87400 73440 1 0 $X=87210 $Y=70480
X955 1 2 70 ICV_16 $T=88320 40800 1 0 $X=88130 $Y=37840
X956 1 2 66 ICV_16 $T=91080 73440 0 0 $X=90890 $Y=73200
X957 1 2 392 ICV_16 $T=95680 40800 1 0 $X=95490 $Y=37840
X958 1 2 84 ICV_16 $T=100280 68000 0 0 $X=100090 $Y=67760
X959 1 2 89 ICV_16 $T=106720 68000 0 0 $X=106530 $Y=67760
X960 1 2 383 ICV_16 $T=119140 40800 0 0 $X=118950 $Y=40560
X961 1 2 103 ICV_16 $T=121900 40800 1 0 $X=121710 $Y=37840
X962 1 2 420 ICV_16 $T=141220 57120 1 0 $X=141030 $Y=54160
X963 1 2 385 ICV_16 $T=142600 46240 1 0 $X=142410 $Y=43280
X964 1 2 130 ICV_16 $T=150880 73440 0 0 $X=150690 $Y=73200
X965 1 2 429 ICV_16 $T=161920 51680 0 0 $X=161730 $Y=51440
X966 1 2 148 ICV_16 $T=181240 46240 1 0 $X=181050 $Y=43280
X967 1 2 154 ICV_16 $T=202400 57120 1 0 $X=202210 $Y=54160
X968 1 2 450 ICV_16 $T=207460 62560 1 0 $X=207270 $Y=59600
X969 1 2 171 ICV_16 $T=208380 40800 1 0 $X=208190 $Y=37840
X970 1 2 154 ICV_16 $T=209760 40800 0 0 $X=209570 $Y=40560
X971 1 2 169 ICV_16 $T=209760 62560 0 0 $X=209570 $Y=62320
X972 1 2 156 ICV_16 $T=210680 35360 0 0 $X=210490 $Y=35120
X973 1 2 6 ICV_16 $T=222180 57120 0 0 $X=221990 $Y=56880
X974 1 2 448 ICV_16 $T=223100 78880 1 0 $X=222910 $Y=75920
X975 1 2 182 ICV_16 $T=231840 57120 0 0 $X=231650 $Y=56880
X976 1 2 165 ICV_16 $T=237820 73440 0 0 $X=237630 $Y=73200
X977 1 2 190 ICV_16 $T=248860 35360 0 0 $X=248670 $Y=35120
X978 1 2 466 ICV_16 $T=251620 51680 0 0 $X=251430 $Y=51440
X979 1 2 478 ICV_16 $T=253000 57120 1 0 $X=252810 $Y=54160
X980 1 2 449 ICV_16 $T=265880 62560 1 0 $X=265690 $Y=59600
X981 1 2 207 ICV_16 $T=273700 40800 0 0 $X=273510 $Y=40560
X982 1 2 501 ICV_16 $T=286580 51680 1 0 $X=286390 $Y=48720
X983 1 2 502 ICV_16 $T=292100 57120 1 0 $X=291910 $Y=54160
X984 1 2 237 ICV_16 $T=308660 46240 1 0 $X=308470 $Y=43280
X985 1 2 342 ICV_16 $T=318780 62560 1 0 $X=318590 $Y=59600
X986 1 2 517 ICV_16 $T=320620 62560 0 0 $X=320430 $Y=62320
X987 1 2 245 ICV_16 $T=322000 68000 0 0 $X=321810 $Y=67760
X988 1 2 525 ICV_16 $T=327520 35360 0 0 $X=327330 $Y=35120
X989 1 2 525 ICV_16 $T=327520 57120 0 0 $X=327330 $Y=56880
X990 1 2 34 2 352 1 sky130_fd_sc_hd__inv_8 $T=32660 73440 1 0 $X=32470 $Y=70480
X991 1 2 28 2 36 1 sky130_fd_sc_hd__inv_8 $T=34500 78880 1 0 $X=34310 $Y=75920
X992 1 2 33 2 353 1 sky130_fd_sc_hd__inv_8 $T=34960 57120 0 0 $X=34770 $Y=56880
X993 1 2 37 2 38 1 sky130_fd_sc_hd__inv_8 $T=39560 40800 1 0 $X=39370 $Y=37840
X994 1 2 43 2 45 1 sky130_fd_sc_hd__inv_8 $T=51520 73440 0 0 $X=51330 $Y=73200
X995 1 2 50 2 56 1 sky130_fd_sc_hd__inv_8 $T=62560 46240 1 0 $X=62370 $Y=43280
X996 1 2 63 2 375 1 sky130_fd_sc_hd__inv_8 $T=74060 35360 0 0 $X=73870 $Y=35120
X997 1 2 85 2 389 1 sky130_fd_sc_hd__inv_8 $T=99820 40800 0 0 $X=99630 $Y=40560
X998 1 2 96 2 399 1 sky130_fd_sc_hd__inv_8 $T=115460 51680 1 0 $X=115270 $Y=48720
X999 1 2 111 2 403 1 sky130_fd_sc_hd__inv_8 $T=133400 46240 1 0 $X=133210 $Y=43280
X1000 1 2 126 2 109 1 sky130_fd_sc_hd__inv_8 $T=149960 35360 0 0 $X=149770 $Y=35120
X1001 1 2 134 2 395 1 sky130_fd_sc_hd__inv_8 $T=161460 62560 1 0 $X=161270 $Y=59600
X1002 1 2 3 2 433 1 sky130_fd_sc_hd__inv_8 $T=166060 46240 0 0 $X=165870 $Y=46000
X1003 1 2 123 2 437 1 sky130_fd_sc_hd__inv_8 $T=166520 40800 1 0 $X=166330 $Y=37840
X1004 1 2 429 2 438 1 sky130_fd_sc_hd__inv_8 $T=168360 62560 1 0 $X=168170 $Y=59600
X1005 1 2 144 2 148 1 sky130_fd_sc_hd__inv_8 $T=175260 35360 0 0 $X=175070 $Y=35120
X1006 1 2 410 2 330 1 sky130_fd_sc_hd__inv_8 $T=179400 51680 1 0 $X=179210 $Y=48720
X1007 1 2 434 2 149 1 sky130_fd_sc_hd__inv_8 $T=183080 62560 0 0 $X=182890 $Y=62320
X1008 1 2 5 2 427 1 sky130_fd_sc_hd__inv_8 $T=185380 68000 0 0 $X=185190 $Y=67760
X1009 1 2 120 2 159 1 sky130_fd_sc_hd__inv_8 $T=211140 73440 0 0 $X=210950 $Y=73200
X1010 1 2 459 2 454 1 sky130_fd_sc_hd__inv_8 $T=214360 51680 0 0 $X=214170 $Y=51440
X1011 1 2 179 2 463 1 sky130_fd_sc_hd__inv_8 $T=220800 35360 0 0 $X=220610 $Y=35120
X1012 1 2 6 2 466 1 sky130_fd_sc_hd__inv_8 $T=222180 62560 1 0 $X=221990 $Y=59600
X1013 1 2 137 2 470 1 sky130_fd_sc_hd__inv_8 $T=239200 68000 0 0 $X=239010 $Y=67760
X1014 1 2 190 2 469 1 sky130_fd_sc_hd__inv_8 $T=245640 40800 1 0 $X=245450 $Y=37840
X1015 1 2 192 2 157 1 sky130_fd_sc_hd__inv_8 $T=245640 62560 1 0 $X=245450 $Y=59600
X1016 1 2 187 2 189 1 sky130_fd_sc_hd__inv_8 $T=245640 78880 1 0 $X=245450 $Y=75920
X1017 1 2 195 2 487 1 sky130_fd_sc_hd__inv_8 $T=260820 40800 0 0 $X=260630 $Y=40560
X1018 1 2 207 2 492 1 sky130_fd_sc_hd__inv_8 $T=273700 46240 1 0 $X=273510 $Y=43280
X1019 1 2 196 2 213 1 sky130_fd_sc_hd__inv_8 $T=273700 73440 1 0 $X=273510 $Y=70480
X1020 1 2 218 2 495 1 sky130_fd_sc_hd__inv_8 $T=278300 57120 0 0 $X=278110 $Y=56880
X1021 1 2 226 2 510 1 sky130_fd_sc_hd__inv_8 $T=301760 51680 1 0 $X=301570 $Y=48720
X1022 1 2 342 2 514 1 sky130_fd_sc_hd__inv_8 $T=315100 68000 1 0 $X=314910 $Y=65040
X1023 1 2 245 2 239 1 sky130_fd_sc_hd__inv_8 $T=320620 78880 1 0 $X=320430 $Y=75920
X1024 1 2 349 346 2 344 1 sky130_fd_sc_hd__nor2_4 $T=32660 62560 1 0 $X=32470 $Y=59600
X1025 1 2 349 348 2 345 1 sky130_fd_sc_hd__nor2_4 $T=34960 51680 0 0 $X=34770 $Y=51440
X1026 1 2 349 350 2 343 1 sky130_fd_sc_hd__nor2_4 $T=34960 62560 0 0 $X=34770 $Y=62320
X1027 1 2 349 347 2 351 1 sky130_fd_sc_hd__nor2_4 $T=36340 51680 1 0 $X=36150 $Y=48720
X1028 1 2 349 355 2 354 1 sky130_fd_sc_hd__nor2_4 $T=40020 68000 1 0 $X=39830 $Y=65040
X1029 1 2 51 371 2 359 1 sky130_fd_sc_hd__nor2_4 $T=63020 51680 0 0 $X=62830 $Y=51440
X1030 1 2 55 60 2 59 1 sky130_fd_sc_hd__nor2_4 $T=66240 35360 0 0 $X=66050 $Y=35120
X1031 1 2 57 372 2 363 1 sky130_fd_sc_hd__nor2_4 $T=66240 62560 1 0 $X=66050 $Y=59600
X1032 1 2 57 61 2 366 1 sky130_fd_sc_hd__nor2_4 $T=67620 62560 0 0 $X=67430 $Y=62320
X1033 1 2 57 65 2 365 1 sky130_fd_sc_hd__nor2_4 $T=72220 68000 0 0 $X=72030 $Y=67760
X1034 1 2 57 71 2 370 1 sky130_fd_sc_hd__nor2_4 $T=77280 62560 1 0 $X=77090 $Y=59600
X1035 1 2 372 385 2 373 1 sky130_fd_sc_hd__nor2_4 $T=81880 51680 0 0 $X=81690 $Y=51440
X1036 1 2 61 385 2 376 1 sky130_fd_sc_hd__nor2_4 $T=81880 57120 0 0 $X=81690 $Y=56880
X1037 1 2 71 385 2 379 1 sky130_fd_sc_hd__nor2_4 $T=91540 57120 1 0 $X=91350 $Y=54160
X1038 1 2 81 391 2 392 1 sky130_fd_sc_hd__nor2_4 $T=93380 51680 1 0 $X=93190 $Y=48720
X1039 1 2 65 84 2 387 1 sky130_fd_sc_hd__nor2_4 $T=95220 68000 0 0 $X=95030 $Y=67760
X1040 1 2 51 394 2 393 1 sky130_fd_sc_hd__nor2_4 $T=101660 57120 0 0 $X=101470 $Y=56880
X1041 1 2 87 86 2 386 1 sky130_fd_sc_hd__nor2_4 $T=104880 73440 0 0 $X=104690 $Y=73200
X1042 1 2 51 396 2 91 1 sky130_fd_sc_hd__nor2_4 $T=105340 46240 1 0 $X=105150 $Y=43280
X1043 1 2 87 98 2 404 1 sky130_fd_sc_hd__nor2_4 $T=115920 73440 1 0 $X=115730 $Y=70480
X1044 1 2 86 106 2 416 1 sky130_fd_sc_hd__nor2_4 $T=127420 73440 0 0 $X=127230 $Y=73200
X1045 1 2 98 106 2 409 1 sky130_fd_sc_hd__nor2_4 $T=133400 78880 1 0 $X=133210 $Y=75920
X1046 1 2 101 422 2 119 1 sky130_fd_sc_hd__nor2_4 $T=138460 40800 1 0 $X=138270 $Y=37840
X1047 1 2 122 385 2 413 1 sky130_fd_sc_hd__nor2_4 $T=142600 51680 1 0 $X=142410 $Y=48720
X1048 1 2 101 421 2 125 1 sky130_fd_sc_hd__nor2_4 $T=146280 40800 1 0 $X=146090 $Y=37840
X1049 1 2 122 414 2 430 1 sky130_fd_sc_hd__nor2_4 $T=149960 57120 0 0 $X=149770 $Y=56880
X1050 1 2 6 334 2 447 1 sky130_fd_sc_hd__nor2_4 $T=189520 57120 1 0 $X=189330 $Y=54160
X1051 1 2 163 452 2 457 1 sky130_fd_sc_hd__nor2_4 $T=203320 46240 0 0 $X=203130 $Y=46000
X1052 1 2 145 170 2 332 1 sky130_fd_sc_hd__nor2_4 $T=203320 73440 0 0 $X=203130 $Y=73200
X1053 1 2 173 461 2 174 1 sky130_fd_sc_hd__nor2_4 $T=219420 40800 1 0 $X=219230 $Y=37840
X1054 1 2 173 473 2 184 1 sky130_fd_sc_hd__nor2_4 $T=230920 40800 1 0 $X=230730 $Y=37840
X1055 1 2 173 468 2 185 1 sky130_fd_sc_hd__nor2_4 $T=231380 40800 0 0 $X=231190 $Y=40560
X1056 1 2 484 482 2 205 1 sky130_fd_sc_hd__nor2_4 $T=259900 46240 1 0 $X=259710 $Y=43280
X1057 1 2 490 491 2 212 1 sky130_fd_sc_hd__nor2_4 $T=268640 40800 0 0 $X=268450 $Y=40560
X1058 1 2 499 501 2 496 1 sky130_fd_sc_hd__nor2_4 $T=287500 51680 0 0 $X=287310 $Y=51440
X1059 1 2 509 511 2 505 1 sky130_fd_sc_hd__nor2_4 $T=297620 57120 0 0 $X=297430 $Y=56880
X1060 1 2 240 516 2 242 1 sky130_fd_sc_hd__nor2_4 $T=310500 78880 1 0 $X=310310 $Y=75920
X1061 1 2 518 517 2 519 1 sky130_fd_sc_hd__nor2_4 $T=315560 62560 0 0 $X=315370 $Y=62320
X1062 1 2 241 522 2 524 1 sky130_fd_sc_hd__nor2_4 $T=315560 73440 0 0 $X=315370 $Y=73200
X1063 1 2 38 329 39 360 2 347 1 sky130_fd_sc_hd__o22a_4 $T=47380 51680 0 0 $X=47190 $Y=51440
X1064 1 2 353 329 39 358 2 348 1 sky130_fd_sc_hd__o22a_4 $T=47840 57120 0 0 $X=47650 $Y=56880
X1065 1 2 36 42 39 361 2 350 1 sky130_fd_sc_hd__o22a_4 $T=49220 68000 1 0 $X=49030 $Y=65040
X1066 1 2 45 42 39 357 2 355 1 sky130_fd_sc_hd__o22a_4 $T=49220 73440 1 0 $X=49030 $Y=70480
X1067 1 2 48 364 38 363 2 360 1 sky130_fd_sc_hd__o22a_4 $T=57040 57120 1 0 $X=56850 $Y=54160
X1068 1 2 48 362 36 366 2 361 1 sky130_fd_sc_hd__o22a_4 $T=58420 68000 1 0 $X=58230 $Y=65040
X1069 1 2 48 369 45 365 2 357 1 sky130_fd_sc_hd__o22a_4 $T=63020 68000 0 0 $X=62830 $Y=67760
X1070 1 2 367 48 353 370 2 358 1 sky130_fd_sc_hd__o22a_4 $T=64400 57120 0 0 $X=64210 $Y=56880
X1071 1 2 56 58 374 368 2 371 1 sky130_fd_sc_hd__o22a_4 $T=65780 73440 1 0 $X=65590 $Y=70480
X1072 1 2 66 58 374 68 2 62 1 sky130_fd_sc_hd__o22a_4 $T=70840 73440 0 0 $X=70650 $Y=73200
X1073 1 2 69 73 56 75 2 368 1 sky130_fd_sc_hd__o22a_4 $T=77280 78880 1 0 $X=77090 $Y=75920
X1074 1 2 364 377 67 373 2 382 1 sky130_fd_sc_hd__o22a_4 $T=78660 46240 0 0 $X=78470 $Y=46000
X1075 1 2 375 383 381 380 2 60 1 sky130_fd_sc_hd__o22a_4 $T=79580 40800 0 0 $X=79390 $Y=40560
X1076 1 2 367 377 375 379 2 380 1 sky130_fd_sc_hd__o22a_4 $T=80040 51680 1 0 $X=79850 $Y=48720
X1077 1 2 67 70 381 382 2 74 1 sky130_fd_sc_hd__o22a_4 $T=80960 40800 1 0 $X=80770 $Y=37840
X1078 1 2 362 377 64 376 2 384 1 sky130_fd_sc_hd__o22a_4 $T=81420 57120 1 0 $X=81230 $Y=54160
X1079 1 2 64 70 381 384 2 76 1 sky130_fd_sc_hd__o22a_4 $T=84640 46240 1 0 $X=84450 $Y=43280
X1080 1 2 69 388 66 386 2 68 1 sky130_fd_sc_hd__o22a_4 $T=87400 78880 1 0 $X=87210 $Y=75920
X1081 1 2 369 377 389 387 2 390 1 sky130_fd_sc_hd__o22a_4 $T=89700 62560 1 0 $X=89510 $Y=59600
X1082 1 2 389 70 381 390 2 391 1 sky130_fd_sc_hd__o22a_4 $T=92000 51680 0 0 $X=91810 $Y=51440
X1083 1 2 90 383 374 397 2 396 1 sky130_fd_sc_hd__o22a_4 $T=105340 51680 1 0 $X=105150 $Y=48720
X1084 1 2 399 383 374 402 2 394 1 sky130_fd_sc_hd__o22a_4 $T=108100 57120 1 0 $X=107910 $Y=54160
X1085 1 2 69 398 90 404 2 397 1 sky130_fd_sc_hd__o22a_4 $T=110860 68000 1 0 $X=110670 $Y=65040
X1086 1 2 94 383 381 400 2 97 1 sky130_fd_sc_hd__o22a_4 $T=114540 40800 1 0 $X=114350 $Y=37840
X1087 1 2 403 383 374 401 2 100 1 sky130_fd_sc_hd__o22a_4 $T=115000 46240 1 0 $X=114810 $Y=43280
X1088 1 2 411 377 403 413 2 401 1 sky130_fd_sc_hd__o22a_4 $T=126960 46240 0 0 $X=126770 $Y=46000
X1089 1 2 398 105 109 409 2 415 1 sky130_fd_sc_hd__o22a_4 $T=128800 68000 0 0 $X=128610 $Y=67760
X1090 1 2 388 105 114 416 2 420 1 sky130_fd_sc_hd__o22a_4 $T=133400 73440 1 0 $X=133210 $Y=70480
X1091 1 2 109 419 115 415 2 421 1 sky130_fd_sc_hd__o22a_4 $T=135700 57120 0 0 $X=135510 $Y=56880
X1092 1 2 114 419 115 420 2 422 1 sky130_fd_sc_hd__o22a_4 $T=137540 62560 1 0 $X=137350 $Y=59600
X1093 1 2 352 423 378 424 2 346 1 sky130_fd_sc_hd__o22a_4 $T=144900 68000 1 0 $X=144710 $Y=65040
X1094 1 2 427 120 99 426 2 423 1 sky130_fd_sc_hd__o22a_4 $T=149040 68000 0 0 $X=148850 $Y=67760
X1095 1 2 72 411 129 430 2 431 1 sky130_fd_sc_hd__o22a_4 $T=151800 62560 0 0 $X=151610 $Y=62320
X1096 1 2 153 156 160 446 2 155 1 sky130_fd_sc_hd__o22a_4 $T=190440 35360 0 0 $X=190250 $Y=35120
X1097 1 2 158 156 160 161 2 164 1 sky130_fd_sc_hd__o22a_4 $T=201020 40800 1 0 $X=200830 $Y=37840
X1098 1 2 454 156 160 455 2 452 1 sky130_fd_sc_hd__o22a_4 $T=202860 51680 1 0 $X=202670 $Y=48720
X1099 1 2 171 156 160 166 2 167 1 sky130_fd_sc_hd__o22a_4 $T=203320 35360 0 0 $X=203130 $Y=35120
X1100 1 2 463 178 175 462 2 461 1 sky130_fd_sc_hd__o22a_4 $T=220340 46240 1 0 $X=220150 $Y=43280
X1101 1 2 469 178 175 471 2 468 1 sky130_fd_sc_hd__o22a_4 $T=230000 51680 1 0 $X=229810 $Y=48720
X1102 1 2 182 178 175 472 2 473 1 sky130_fd_sc_hd__o22a_4 $T=231380 46240 0 0 $X=231190 $Y=46000
X1103 1 2 356 2 349 1 sky130_fd_sc_hd__buf_1 $T=49220 57120 1 0 $X=49030 $Y=54160
X1104 1 2 356 2 44 1 sky130_fd_sc_hd__buf_1 $T=49220 78880 1 0 $X=49030 $Y=75920
X1105 1 2 356 2 51 1 sky130_fd_sc_hd__buf_1 $T=60720 51680 1 0 $X=60530 $Y=48720
X1106 1 2 49 2 329 1 sky130_fd_sc_hd__buf_1 $T=61180 62560 1 0 $X=60990 $Y=59600
X1107 1 2 53 2 39 1 sky130_fd_sc_hd__buf_1 $T=63020 62560 0 0 $X=62830 $Y=62320
X1108 1 2 49 2 42 1 sky130_fd_sc_hd__buf_1 $T=63020 73440 0 0 $X=62830 $Y=73200
X1109 1 2 49 2 58 1 sky130_fd_sc_hd__buf_1 $T=67160 78880 1 0 $X=66970 $Y=75920
X1110 1 2 356 2 55 1 sky130_fd_sc_hd__buf_1 $T=77280 46240 1 0 $X=77090 $Y=43280
X1111 1 2 53 2 374 1 sky130_fd_sc_hd__buf_1 $T=77280 57120 1 0 $X=77090 $Y=54160
X1112 1 2 69 2 48 1 sky130_fd_sc_hd__buf_1 $T=77280 73440 1 0 $X=77090 $Y=70480
X1113 1 2 72 2 57 1 sky130_fd_sc_hd__buf_1 $T=80040 68000 0 0 $X=79850 $Y=67760
X1114 1 2 356 2 81 1 sky130_fd_sc_hd__buf_1 $T=97980 62560 0 0 $X=97790 $Y=62320
X1115 1 2 395 2 356 1 sky130_fd_sc_hd__buf_1 $T=103040 62560 0 0 $X=102850 $Y=62320
X1116 1 2 49 2 383 1 sky130_fd_sc_hd__buf_1 $T=105340 62560 1 0 $X=105150 $Y=59600
X1117 1 2 89 2 70 1 sky130_fd_sc_hd__buf_1 $T=106720 73440 1 0 $X=106530 $Y=70480
X1118 1 2 95 2 78 1 sky130_fd_sc_hd__buf_1 $T=112700 73440 0 0 $X=112510 $Y=73200
X1119 1 2 99 2 381 1 sky130_fd_sc_hd__buf_1 $T=115920 62560 1 0 $X=115730 $Y=59600
X1120 1 2 395 2 101 1 sky130_fd_sc_hd__buf_1 $T=119140 57120 0 0 $X=118950 $Y=56880
X1121 1 2 405 2 84 1 sky130_fd_sc_hd__buf_1 $T=119140 68000 0 0 $X=118950 $Y=67760
X1122 1 2 408 2 69 1 sky130_fd_sc_hd__buf_1 $T=120980 68000 1 0 $X=120790 $Y=65040
X1123 1 2 105 2 377 1 sky130_fd_sc_hd__buf_1 $T=122820 62560 0 0 $X=122630 $Y=62320
X1124 1 2 405 2 106 1 sky130_fd_sc_hd__buf_1 $T=126500 73440 1 0 $X=126310 $Y=70480
X1125 1 2 108 2 105 1 sky130_fd_sc_hd__buf_1 $T=126960 78880 1 0 $X=126770 $Y=75920
X1126 1 2 414 2 87 1 sky130_fd_sc_hd__buf_1 $T=133400 62560 1 0 $X=133210 $Y=59600
X1127 1 2 99 2 115 1 sky130_fd_sc_hd__buf_1 $T=135240 73440 0 0 $X=135050 $Y=73200
X1128 1 2 405 2 385 1 sky130_fd_sc_hd__buf_1 $T=137080 51680 1 0 $X=136890 $Y=48720
X1129 1 2 414 2 72 1 sky130_fd_sc_hd__buf_1 $T=140760 62560 0 0 $X=140570 $Y=62320
X1130 1 2 425 2 405 1 sky130_fd_sc_hd__buf_1 $T=147200 51680 0 0 $X=147010 $Y=51440
X1131 1 2 130 2 131 1 sky130_fd_sc_hd__buf_1 $T=150880 78880 1 0 $X=150690 $Y=75920
X1132 1 2 428 2 414 1 sky130_fd_sc_hd__buf_1 $T=151800 51680 0 0 $X=151610 $Y=51440
X1133 1 2 128 2 99 1 sky130_fd_sc_hd__buf_1 $T=155020 73440 1 0 $X=154830 $Y=70480
X1134 1 2 136 2 410 1 sky130_fd_sc_hd__buf_1 $T=161460 73440 1 0 $X=161270 $Y=70480
X1135 1 2 429 2 412 1 sky130_fd_sc_hd__buf_1 $T=161920 57120 1 0 $X=161730 $Y=54160
X1136 1 2 132 2 378 1 sky130_fd_sc_hd__buf_1 $T=163300 46240 1 0 $X=163110 $Y=43280
X1137 1 2 436 2 429 1 sky130_fd_sc_hd__buf_1 $T=164680 57120 0 0 $X=164490 $Y=56880
X1138 1 2 438 2 49 1 sky130_fd_sc_hd__buf_1 $T=168820 62560 0 0 $X=168630 $Y=62320
X1139 1 2 132 2 95 1 sky130_fd_sc_hd__buf_1 $T=169280 46240 1 0 $X=169090 $Y=43280
X1140 1 2 412 2 145 1 sky130_fd_sc_hd__buf_1 $T=176180 62560 1 0 $X=175990 $Y=59600
X1141 1 2 438 2 89 1 sky130_fd_sc_hd__buf_1 $T=189520 73440 1 0 $X=189330 $Y=70480
X1142 1 2 89 2 419 1 sky130_fd_sc_hd__buf_1 $T=193660 73440 1 0 $X=193470 $Y=70480
X1143 1 2 453 2 434 1 sky130_fd_sc_hd__buf_1 $T=196420 68000 1 0 $X=196230 $Y=65040
X1144 1 2 450 2 6 1 sky130_fd_sc_hd__buf_1 $T=201480 62560 1 0 $X=201290 $Y=59600
X1145 1 2 7 2 5 1 sky130_fd_sc_hd__buf_1 $T=207000 78880 1 0 $X=206810 $Y=75920
X1146 1 2 128 2 53 1 sky130_fd_sc_hd__buf_1 $T=231380 68000 0 0 $X=231190 $Y=67760
X1147 1 2 165 2 449 1 sky130_fd_sc_hd__buf_1 $T=232760 78880 1 0 $X=232570 $Y=75920
X1148 1 2 165 2 177 1 sky130_fd_sc_hd__buf_1 $T=237820 78880 1 0 $X=237630 $Y=75920
X1149 1 2 192 2 169 1 sky130_fd_sc_hd__buf_1 $T=252080 57120 0 0 $X=251890 $Y=56880
X1150 1 2 486 2 187 1 sky130_fd_sc_hd__buf_1 $T=262660 73440 0 0 $X=262470 $Y=73200
X1151 1 2 169 2 214 1 sky130_fd_sc_hd__buf_1 $T=270020 73440 0 0 $X=269830 $Y=73200
X1152 1 2 196 2 198 1 sky130_fd_sc_hd__buf_1 $T=274620 68000 0 0 $X=274430 $Y=67760
X1153 1 2 206 2 215 1 sky130_fd_sc_hd__buf_1 $T=275540 78880 1 0 $X=275350 $Y=75920
X1154 1 2 216 2 483 1 sky130_fd_sc_hd__buf_1 $T=280600 62560 0 0 $X=280410 $Y=62320
X1155 1 2 216 2 188 1 sky130_fd_sc_hd__buf_1 $T=281060 68000 1 0 $X=280870 $Y=65040
X1156 1 2 202 2 498 1 sky130_fd_sc_hd__buf_1 $T=281980 73440 1 0 $X=281790 $Y=70480
X1157 1 2 216 2 221 1 sky130_fd_sc_hd__buf_1 $T=287960 68000 0 0 $X=287770 $Y=67760
X1158 1 2 437 433 410 2 141 1 sky130_fd_sc_hd__o21a_4 $T=170200 51680 1 0 $X=170010 $Y=48720
X1159 1 2 148 410 385 2 439 1 sky130_fd_sc_hd__o21a_4 $T=175260 46240 0 0 $X=175070 $Y=46000
X1160 1 2 104 153 154 2 446 1 sky130_fd_sc_hd__o21a_4 $T=189520 40800 1 0 $X=189330 $Y=37840
X1161 1 2 102 158 154 2 161 1 sky130_fd_sc_hd__o21a_4 $T=199180 46240 1 0 $X=198990 $Y=43280
X1162 1 2 82 171 154 2 166 1 sky130_fd_sc_hd__o21a_4 $T=203320 40800 0 0 $X=203130 $Y=40560
X1163 1 2 107 454 154 2 455 1 sky130_fd_sc_hd__o21a_4 $T=203320 51680 0 0 $X=203130 $Y=51440
X1164 1 2 159 5 4 2 458 1 sky130_fd_sc_hd__o21a_4 $T=207000 73440 1 0 $X=206810 $Y=70480
X1165 1 2 139 463 180 2 462 1 sky130_fd_sc_hd__o21a_4 $T=220800 51680 1 0 $X=220610 $Y=48720
X1166 1 2 466 465 451 2 467 1 sky130_fd_sc_hd__o21a_4 $T=226320 73440 1 0 $X=226130 $Y=70480
X1167 1 2 181 469 180 2 471 1 sky130_fd_sc_hd__o21a_4 $T=231380 51680 0 0 $X=231190 $Y=51440
X1168 1 2 146 182 180 2 472 1 sky130_fd_sc_hd__o21a_4 $T=231840 57120 1 0 $X=231650 $Y=54160
X1169 1 2 466 474 476 2 475 1 sky130_fd_sc_hd__o21a_4 $T=242880 57120 0 0 $X=242690 $Y=56880
X1170 1 2 466 477 479 2 478 1 sky130_fd_sc_hd__o21a_4 $T=247940 62560 0 0 $X=247750 $Y=62320
X1171 1 2 364 ICV_22 $T=55660 51680 1 0 $X=55470 $Y=48720
X1172 1 2 8 ICV_22 $T=118220 35360 0 0 $X=118030 $Y=35120
X1173 1 2 86 ICV_22 $T=124200 73440 0 0 $X=124010 $Y=73200
X1174 1 2 414 ICV_22 $T=126040 62560 0 0 $X=125850 $Y=62320
X1175 1 2 116 ICV_22 $T=137540 78880 1 0 $X=137350 $Y=75920
X1176 1 2 113 ICV_22 $T=148580 51680 0 0 $X=148390 $Y=51440
X1177 1 2 89 ICV_22 $T=186760 73440 0 0 $X=186570 $Y=73200
X1178 1 2 438 ICV_22 $T=202400 62560 0 0 $X=202210 $Y=62320
X1179 1 2 8 ICV_22 $T=207460 46240 0 0 $X=207270 $Y=46000
X1180 1 2 338 ICV_22 $T=208840 57120 1 0 $X=208650 $Y=54160
X1181 1 2 8 ICV_22 $T=234140 35360 0 0 $X=233950 $Y=35120
X1182 1 2 8 ICV_22 $T=237820 46240 0 0 $X=237630 $Y=46000
X1183 1 2 188 ICV_22 $T=244720 51680 1 0 $X=244530 $Y=48720
X1184 1 2 198 ICV_22 $T=249780 62560 1 0 $X=249590 $Y=59600
X1185 1 2 225 ICV_22 $T=291640 51680 0 0 $X=291450 $Y=51440
X1186 1 2 227 ICV_22 $T=293020 78880 1 0 $X=292830 $Y=75920
X1187 1 2 523 ICV_22 $T=320160 46240 0 0 $X=319970 $Y=46000
X1188 1 2 521 ICV_22 $T=320620 35360 0 0 $X=320430 $Y=35120
X1189 1 2 525 ICV_22 $T=328900 40800 1 0 $X=328710 $Y=37840
X1190 1 2 ICV_26 $T=5520 35360 0 0 $X=5330 $Y=35120
X1191 1 2 ICV_26 $T=5520 40800 0 0 $X=5330 $Y=40560
X1192 1 2 ICV_26 $T=5520 46240 0 0 $X=5330 $Y=46000
X1193 1 2 ICV_26 $T=5520 51680 0 0 $X=5330 $Y=51440
X1194 1 2 ICV_26 $T=5520 57120 0 0 $X=5330 $Y=56880
X1195 1 2 ICV_26 $T=5520 62560 0 0 $X=5330 $Y=62320
X1196 1 2 ICV_26 $T=5520 68000 0 0 $X=5330 $Y=67760
X1197 1 2 ICV_26 $T=5520 73440 0 0 $X=5330 $Y=73200
X1198 1 2 ICV_26 $T=350520 35360 1 180 $X=348950 $Y=35120
X1199 1 2 ICV_26 $T=350520 40800 1 180 $X=348950 $Y=40560
X1200 1 2 ICV_26 $T=350520 46240 1 180 $X=348950 $Y=46000
X1201 1 2 ICV_26 $T=350520 51680 1 180 $X=348950 $Y=51440
X1202 1 2 ICV_26 $T=350520 57120 1 180 $X=348950 $Y=56880
X1203 1 2 ICV_26 $T=350520 62560 1 180 $X=348950 $Y=62320
X1204 1 2 ICV_26 $T=350520 68000 1 180 $X=348950 $Y=67760
X1205 1 2 ICV_26 $T=350520 73440 1 180 $X=348950 $Y=73200
X1206 1 2 36 361 ICV_27 $T=50140 62560 0 0 $X=49950 $Y=62320
X1207 1 2 374 66 ICV_27 $T=70840 78880 1 0 $X=70650 $Y=75920
X1208 1 2 380 356 ICV_27 $T=74520 40800 0 0 $X=74330 $Y=40560
X1209 1 2 378 53 ICV_27 $T=76820 51680 0 0 $X=76630 $Y=51440
X1210 1 2 367 383 ICV_27 $T=80040 46240 1 0 $X=79850 $Y=43280
X1211 1 2 381 390 ICV_27 $T=96600 57120 1 0 $X=96410 $Y=54160
X1212 1 2 90 397 ICV_27 $T=107180 46240 0 0 $X=106990 $Y=46000
X1213 1 2 90 404 ICV_27 $T=112700 62560 0 0 $X=112510 $Y=62320
X1214 1 2 403 377 ICV_27 $T=126960 46240 1 0 $X=126770 $Y=43280
X1215 1 2 109 105 ICV_27 $T=126960 68000 1 0 $X=126770 $Y=65040
X1216 1 2 418 417 ICV_27 $T=133400 40800 1 0 $X=133210 $Y=37840
X1217 1 2 116 121 ICV_27 $T=140760 73440 0 0 $X=140570 $Y=73200
X1218 1 2 132 122 ICV_27 $T=153180 46240 1 0 $X=152990 $Y=43280
X1219 1 2 142 145 ICV_27 $T=173420 78880 1 0 $X=173230 $Y=75920
X1220 1 2 157 118 ICV_27 $T=195040 73440 0 0 $X=194850 $Y=73200
X1221 1 2 165 168 ICV_27 $T=202400 78880 1 0 $X=202210 $Y=75920
X1222 1 2 450 332 ICV_27 $T=203320 57120 0 0 $X=203130 $Y=56880
X1223 1 2 82 455 ICV_27 $T=205620 46240 1 0 $X=205430 $Y=43280
X1224 1 2 8 467 ICV_27 $T=224940 62560 0 0 $X=224750 $Y=62320
X1225 1 2 195 200 ICV_27 $T=251160 40800 0 0 $X=250970 $Y=40560
X1226 1 2 196 209 ICV_27 $T=264960 73440 0 0 $X=264770 $Y=73200
X1227 1 2 206 217 ICV_27 $T=275540 73440 0 0 $X=275350 $Y=73200
X1228 1 2 210 216 ICV_27 $T=290260 68000 0 0 $X=290070 $Y=67760
X1229 1 2 243 244 ICV_27 $T=315560 78880 1 0 $X=315370 $Y=75920
X1230 1 2 240 516 ICV_27 $T=318320 73440 1 0 $X=318130 $Y=70480
X1231 1 2 38 ICV_28 $T=58880 51680 0 0 $X=58690 $Y=51440
X1232 1 2 374 ICV_28 $T=73140 73440 1 0 $X=72950 $Y=70480
X1233 1 2 381 ICV_28 $T=86940 40800 0 0 $X=86750 $Y=40560
X1234 1 2 372 ICV_28 $T=86940 51680 0 0 $X=86750 $Y=51440
X1235 1 2 374 ICV_28 $T=115000 40800 0 0 $X=114810 $Y=40560
X1236 1 2 95 ICV_28 $T=115000 73440 0 0 $X=114810 $Y=73200
X1237 1 2 95 ICV_28 $T=129260 62560 1 0 $X=129070 $Y=59600
X1238 1 2 114 ICV_28 $T=143060 57120 0 0 $X=142870 $Y=56880
X1239 1 2 414 ICV_28 $T=143060 62560 0 0 $X=142870 $Y=62320
X1240 1 2 433 ICV_28 $T=171120 46240 0 0 $X=170930 $Y=46000
X1241 1 2 438 ICV_28 $T=171120 62560 0 0 $X=170930 $Y=62320
X1242 1 2 102 ICV_28 $T=199180 40800 0 0 $X=198990 $Y=40560
X1243 1 2 120 ICV_28 $T=199180 68000 0 0 $X=198990 $Y=67760
X1244 1 2 196 ICV_28 $T=255300 73440 0 0 $X=255110 $Y=73200
X1245 1 2 509 ICV_28 $T=297620 62560 1 0 $X=297430 $Y=59600
X1246 1 2 525 ICV_28 $T=325680 40800 1 0 $X=325490 $Y=37840
X1247 1 2 521 ICV_28 $T=325680 46240 1 0 $X=325490 $Y=43280
X1248 1 2 7 ICV_28 $T=339480 46240 0 0 $X=339290 $Y=46000
X1249 1 2 ICV_29 $T=10580 40800 1 0 $X=10390 $Y=37840
X1250 1 2 ICV_29 $T=10580 62560 1 0 $X=10390 $Y=59600
X1251 1 2 ICV_29 $T=10580 73440 1 0 $X=10390 $Y=70480
X1252 1 2 ICV_29 $T=10580 78880 1 0 $X=10390 $Y=75920
X1253 1 2 ICV_29 $T=18400 57120 0 0 $X=18210 $Y=56880
X1254 1 2 ICV_29 $T=23000 73440 0 0 $X=22810 $Y=73200
X1255 1 2 ICV_29 $T=38640 78880 1 0 $X=38450 $Y=75920
X1256 1 2 ICV_29 $T=51060 40800 0 0 $X=50870 $Y=40560
X1257 1 2 ICV_29 $T=51060 46240 0 0 $X=50870 $Y=46000
X1258 1 2 ICV_29 $T=93840 78880 1 0 $X=93650 $Y=75920
X1259 1 2 ICV_29 $T=94760 46240 1 0 $X=94570 $Y=43280
X1260 1 2 ICV_29 $T=106720 62560 1 0 $X=106530 $Y=59600
X1261 1 2 ICV_29 $T=150420 40800 1 0 $X=150230 $Y=37840
X1262 1 2 ICV_29 $T=162840 73440 1 0 $X=162650 $Y=70480
X1263 1 2 ICV_29 $T=178020 40800 1 0 $X=177830 $Y=37840
X1264 1 2 ICV_29 $T=192740 57120 0 0 $X=192550 $Y=56880
X1265 1 2 ICV_29 $T=235060 40800 1 0 $X=234870 $Y=37840
X1266 1 2 ICV_29 $T=241040 40800 0 0 $X=240850 $Y=40560
X1267 1 2 ICV_29 $T=249780 40800 1 0 $X=249590 $Y=37840
X1268 1 2 ICV_29 $T=267720 62560 0 0 $X=267530 $Y=62320
X1269 1 2 ICV_29 $T=286580 73440 0 0 $X=286390 $Y=73200
X1270 1 2 ICV_29 $T=305900 51680 1 0 $X=305710 $Y=48720
X1271 1 2 ICV_29 $T=319240 68000 1 0 $X=319050 $Y=65040
X1272 1 2 ICV_29 $T=332580 62560 0 0 $X=332390 $Y=62320
X1273 1 2 ICV_29 $T=339940 68000 1 0 $X=339750 $Y=65040
X1274 1 2 372 378 2 364 1 sky130_fd_sc_hd__or2_4 $T=72680 51680 0 0 $X=72490 $Y=51440
X1275 1 2 61 378 2 362 1 sky130_fd_sc_hd__or2_4 $T=74520 57120 0 0 $X=74330 $Y=56880
X1276 1 2 65 378 2 369 1 sky130_fd_sc_hd__or2_4 $T=77280 62560 0 0 $X=77090 $Y=62320
X1277 1 2 77 375 2 82 1 sky130_fd_sc_hd__or2_4 $T=91080 46240 0 0 $X=90890 $Y=46000
X1278 1 2 77 67 2 79 1 sky130_fd_sc_hd__or2_4 $T=91080 57120 0 0 $X=90890 $Y=56880
X1279 1 2 77 64 2 80 1 sky130_fd_sc_hd__or2_4 $T=91080 62560 0 0 $X=90890 $Y=62320
X1280 1 2 71 78 2 367 1 sky130_fd_sc_hd__or2_4 $T=91080 68000 1 0 $X=90890 $Y=65040
X1281 1 2 77 389 2 83 1 sky130_fd_sc_hd__or2_4 $T=93840 73440 1 0 $X=93650 $Y=70480
X1282 1 2 92 90 2 93 1 sky130_fd_sc_hd__or2_4 $T=109020 78880 1 0 $X=108830 $Y=75920
X1283 1 2 86 78 2 388 1 sky130_fd_sc_hd__or2_4 $T=115920 78880 1 0 $X=115730 $Y=75920
X1284 1 2 92 94 2 102 1 sky130_fd_sc_hd__or2_4 $T=119140 46240 0 0 $X=118950 $Y=46000
X1285 1 2 92 399 2 104 1 sky130_fd_sc_hd__or2_4 $T=119140 51680 0 0 $X=118950 $Y=51440
X1286 1 2 98 78 2 398 1 sky130_fd_sc_hd__or2_4 $T=119140 73440 0 0 $X=118950 $Y=73200
X1287 1 2 92 403 2 107 1 sky130_fd_sc_hd__or2_4 $T=123280 51680 1 0 $X=123090 $Y=48720
X1288 1 2 410 87 2 407 1 sky130_fd_sc_hd__or2_4 $T=125120 62560 1 0 $X=124930 $Y=59600
X1289 1 2 414 412 2 408 1 sky130_fd_sc_hd__or2_4 $T=129260 62560 0 0 $X=129070 $Y=62320
X1290 1 2 405 113 2 418 1 sky130_fd_sc_hd__or2_4 $T=137080 46240 0 0 $X=136890 $Y=46000
X1291 1 2 3 123 2 428 1 sky130_fd_sc_hd__or2_4 $T=149040 46240 0 0 $X=148850 $Y=46000
X1292 1 2 425 429 2 108 1 sky130_fd_sc_hd__or2_4 $T=151800 57120 1 0 $X=151610 $Y=54160
X1293 1 2 122 132 2 411 1 sky130_fd_sc_hd__or2_4 $T=153180 51680 1 0 $X=152990 $Y=48720
X1294 1 2 433 123 2 425 1 sky130_fd_sc_hd__or2_4 $T=158700 46240 0 0 $X=158510 $Y=46000
X1295 1 2 431 99 2 435 1 sky130_fd_sc_hd__or2_4 $T=159160 68000 0 0 $X=158970 $Y=67760
X1296 1 2 120 7 2 436 1 sky130_fd_sc_hd__or2_4 $T=161920 62560 0 0 $X=161730 $Y=62320
X1297 1 2 137 352 2 139 1 sky130_fd_sc_hd__or2_4 $T=164220 68000 1 0 $X=164030 $Y=65040
X1298 1 2 137 353 2 146 1 sky130_fd_sc_hd__or2_4 $T=175260 62560 0 0 $X=175070 $Y=62320
X1299 1 2 149 395 2 450 1 sky130_fd_sc_hd__or2_4 $T=189520 68000 1 0 $X=189330 $Y=65040
X1300 1 2 157 159 2 453 1 sky130_fd_sc_hd__or2_4 $T=195040 68000 0 0 $X=194850 $Y=67760
X1301 1 2 456 450 2 172 1 sky130_fd_sc_hd__or2_4 $T=205620 68000 1 0 $X=205430 $Y=65040
X1302 1 2 474 202 2 204 1 sky130_fd_sc_hd__or2_4 $T=256220 78880 1 0 $X=256030 $Y=75920
X1303 1 2 210 211 2 489 1 sky130_fd_sc_hd__or2_4 $T=264960 68000 1 0 $X=264770 $Y=65040
X1304 1 2 210 187 2 494 1 sky130_fd_sc_hd__or2_4 $T=267720 68000 0 0 $X=267530 $Y=67760
X1305 1 2 210 222 2 500 1 sky130_fd_sc_hd__or2_4 $T=287040 73440 1 0 $X=286850 $Y=70480
X1306 1 2 228 210 2 512 1 sky130_fd_sc_hd__or2_4 $T=297620 73440 0 0 $X=297430 $Y=73200
X1307 1 2 434 432 2 424 1 sky130_fd_sc_hd__and2_4 $T=157780 57120 0 0 $X=157590 $Y=56880
X1308 1 2 169 438 2 456 1 sky130_fd_sc_hd__and2_4 $T=205620 62560 0 0 $X=205430 $Y=62320
X1309 1 2 177 448 2 465 1 sky130_fd_sc_hd__and2_4 $T=223100 73440 0 0 $X=222910 $Y=73200
X1310 1 2 470 183 2 464 1 sky130_fd_sc_hd__and2_4 $T=231380 73440 0 0 $X=231190 $Y=73200
X1311 1 2 115 188 2 476 1 sky130_fd_sc_hd__and2_4 $T=246100 57120 1 0 $X=245910 $Y=54160
X1312 1 2 470 191 2 474 1 sky130_fd_sc_hd__and2_4 $T=247020 68000 0 0 $X=246830 $Y=67760
X1313 1 2 466 474 2 480 1 sky130_fd_sc_hd__and2_4 $T=247480 51680 0 0 $X=247290 $Y=51440
X1314 1 2 194 470 2 477 1 sky130_fd_sc_hd__and2_4 $T=250700 73440 1 0 $X=250510 $Y=70480
X1315 1 2 196 193 2 201 1 sky130_fd_sc_hd__and2_4 $T=251160 73440 0 0 $X=250970 $Y=73200
X1316 1 2 195 200 2 481 1 sky130_fd_sc_hd__and2_4 $T=253000 46240 1 0 $X=252810 $Y=43280
X1317 1 2 207 208 2 488 1 sky130_fd_sc_hd__and2_4 $T=263120 51680 0 0 $X=262930 $Y=51440
X1318 1 2 226 225 2 508 1 sky130_fd_sc_hd__and2_4 $T=294860 51680 0 0 $X=294670 $Y=51440
X1319 1 2 342 230 2 513 1 sky130_fd_sc_hd__and2_4 $T=301760 73440 1 0 $X=301570 $Y=70480
X1320 1 2 87 113 120 2 426 1 sky130_fd_sc_hd__nor3_4 $T=142600 73440 1 0 $X=142410 $Y=70480
X1321 1 2 6 464 458 2 460 1 sky130_fd_sc_hd__nor3_4 $T=217580 73440 1 0 $X=217390 $Y=70480
X1322 1 2 483 481 485 2 484 1 sky130_fd_sc_hd__nor3_4 $T=261280 46240 0 0 $X=261090 $Y=46000
X1323 1 2 483 488 493 2 490 1 sky130_fd_sc_hd__nor3_4 $T=273700 51680 1 0 $X=273510 $Y=48720
X1324 1 2 53 191 495 2 497 1 sky130_fd_sc_hd__nor3_4 $T=276460 62560 1 0 $X=276270 $Y=59600
X1325 1 2 221 497 502 2 499 1 sky130_fd_sc_hd__nor3_4 $T=286120 62560 1 0 $X=285930 $Y=59600
X1326 1 2 221 508 506 2 509 1 sky130_fd_sc_hd__nor3_4 $T=301760 57120 1 0 $X=301570 $Y=54160
X1327 1 2 221 513 507 2 518 1 sky130_fd_sc_hd__nor3_4 $T=302220 68000 0 0 $X=302030 $Y=67760
X1328 1 2 441 443 329 143 2 1 sky130_fd_sc_hd__a21oi_4 $T=174340 46240 1 0 $X=174150 $Y=43280
X1329 1 2 440 434 442 147 2 1 sky130_fd_sc_hd__a21oi_4 $T=175720 73440 1 0 $X=175530 $Y=70480
X1330 1 2 489 449 487 485 2 1 sky130_fd_sc_hd__a21oi_4 $T=265880 57120 0 0 $X=265690 $Y=56880
X1331 1 2 494 449 492 493 2 1 sky130_fd_sc_hd__a21oi_4 $T=270020 51680 0 0 $X=269830 $Y=51440
X1332 1 2 500 177 495 502 2 1 sky130_fd_sc_hd__a21oi_4 $T=287500 62560 0 0 $X=287310 $Y=62320
X1333 1 2 512 177 510 506 2 1 sky130_fd_sc_hd__a21oi_4 $T=300840 62560 0 0 $X=300650 $Y=62320
X1334 1 2 229 449 231 233 2 1 sky130_fd_sc_hd__a21oi_4 $T=301760 78880 1 0 $X=301570 $Y=75920
X1335 1 2 236 177 514 507 2 1 sky130_fd_sc_hd__a21oi_4 $T=307740 73440 1 0 $X=307550 $Y=70480
X1336 1 29 7 ICV_36 $T=29900 35360 0 0 $X=29710 $Y=35120
X1337 1 348 349 ICV_36 $T=29900 51680 0 0 $X=29710 $Y=51440
X1338 1 49 367 ICV_36 $T=57960 57120 0 0 $X=57770 $Y=56880
X1339 1 64 67 ICV_36 $T=72220 51680 1 0 $X=72030 $Y=48720
X1340 1 376 61 ICV_36 $T=72220 57120 1 0 $X=72030 $Y=54160
X1341 1 377 77 ICV_36 $T=86020 46240 0 0 $X=85830 $Y=46000
X1342 1 98 87 ICV_36 $T=114080 68000 0 0 $X=113890 $Y=67760
X1343 1 410 72 ICV_36 $T=128340 57120 1 0 $X=128150 $Y=54160
X1344 1 421 101 ICV_36 $T=142140 35360 0 0 $X=141950 $Y=35120
X1345 1 439 53 ICV_36 $T=170200 51680 0 0 $X=170010 $Y=51440
X1346 1 440 442 ICV_36 $T=170200 68000 0 0 $X=170010 $Y=67760
X1347 1 419 129 ICV_36 $T=170200 73440 0 0 $X=170010 $Y=73200
X1348 1 127 4 ICV_36 $T=184460 78880 1 0 $X=184270 $Y=75920
X1349 1 160 163 ICV_36 $T=198260 46240 0 0 $X=198070 $Y=46000
X1350 1 454 107 ICV_36 $T=198260 51680 0 0 $X=198070 $Y=51440
X1351 1 453 6 ICV_36 $T=198260 62560 0 0 $X=198070 $Y=62320
X1352 1 468 173 ICV_36 $T=226320 40800 0 0 $X=226130 $Y=40560
X1353 1 469 175 ICV_36 $T=226320 46240 0 0 $X=226130 $Y=46000
X1354 1 181 146 ICV_36 $T=226320 51680 0 0 $X=226130 $Y=51440
X1355 1 203 188 ICV_36 $T=268640 46240 1 0 $X=268450 $Y=43280
X1356 1 449 231 ICV_36 $T=296700 73440 1 0 $X=296510 $Y=70480
X1357 1 239 483 ICV_36 $T=310500 68000 0 0 $X=310310 $Y=67760
X1358 1 2 410 95 72 412 2 406 1 sky130_fd_sc_hd__or4_4 $T=127420 57120 0 0 $X=127230 $Y=56880
X1359 1 2 113 95 405 412 2 417 1 sky130_fd_sc_hd__or4_4 $T=134780 51680 0 0 $X=134590 $Y=51440
X1360 1 2 116 118 117 121 2 372 1 sky130_fd_sc_hd__or4_4 $T=140760 78880 1 0 $X=140570 $Y=75920
X1361 1 2 412 128 113 72 2 432 1 sky130_fd_sc_hd__or4_4 $T=149960 62560 1 0 $X=149770 $Y=59600
X1362 1 2 196 209 206 169 2 486 1 sky130_fd_sc_hd__or4_4 $T=263120 78880 1 0 $X=262930 $Y=75920
X1363 1 2 118 419 140 2 451 1 sky130_fd_sc_hd__and3_4 $T=189980 73440 0 0 $X=189790 $Y=73200
X1364 1 2 120 117 449 2 331 1 sky130_fd_sc_hd__and3_4 $T=199180 73440 1 0 $X=198990 $Y=70480
X1365 1 2 219 194 215 2 220 1 sky130_fd_sc_hd__and3_4 $T=280600 78880 1 0 $X=280410 $Y=75920
X1366 1 2 439 445 53 2 443 1 sky130_fd_sc_hd__or3_4 $T=175260 51680 0 0 $X=175070 $Y=51440
X1367 1 2 134 434 123 329 2 135 1 sky130_fd_sc_hd__and4_4 $T=161460 51680 1 0 $X=161270 $Y=48720
X1368 1 2 437 3 330 378 2 445 1 sky130_fd_sc_hd__and4_4 $T=175260 40800 0 0 $X=175070 $Y=40560
X1369 1 2 406 407 96 2 402 1 sky130_fd_sc_hd__a21boi_4 $T=120520 57120 1 0 $X=120330 $Y=54160
X1370 1 2 417 418 110 2 400 1 sky130_fd_sc_hd__a21boi_4 $T=131560 40800 0 0 $X=131370 $Y=40560
X1371 1 2 504 503 2 1 sky130_fd_sc_hd__clkbuf_1 $T=293940 40800 0 0 $X=293750 $Y=40560
X1372 1 2 237 515 2 1 sky130_fd_sc_hd__clkbuf_1 $T=307280 40800 0 0 $X=307090 $Y=40560
X1373 1 2 520 521 2 1 sky130_fd_sc_hd__clkbuf_1 $T=310960 46240 0 0 $X=310770 $Y=46000
X1374 1 2 504 238 2 1 sky130_fd_sc_hd__clkbuf_1 $T=319240 35360 0 0 $X=319050 $Y=35120
X1375 1 2 520 525 2 1 sky130_fd_sc_hd__clkbuf_1 $T=337180 46240 0 0 $X=336990 $Y=46000
X1376 1 2 503 2 551 1 sky130_fd_sc_hd__clkbuf_4 $T=303140 40800 1 0 $X=302950 $Y=37840
X1377 1 2 503 2 552 1 sky130_fd_sc_hd__clkbuf_4 $T=303140 40800 0 0 $X=302950 $Y=40560
X1378 1 2 238 2 553 1 sky130_fd_sc_hd__clkbuf_4 $T=309580 40800 0 0 $X=309390 $Y=40560
X1379 1 2 515 2 523 1 sky130_fd_sc_hd__clkbuf_4 $T=315560 35360 0 0 $X=315370 $Y=35120
X1380 1 2 521 2 554 1 sky130_fd_sc_hd__clkbuf_4 $T=315560 46240 1 0 $X=315370 $Y=43280
X1381 1 2 521 2 555 1 sky130_fd_sc_hd__clkbuf_4 $T=315560 51680 1 0 $X=315370 $Y=48720
X1382 1 2 521 2 556 1 sky130_fd_sc_hd__clkbuf_4 $T=317400 40800 0 0 $X=317210 $Y=40560
X1383 1 2 521 2 557 1 sky130_fd_sc_hd__clkbuf_4 $T=317400 46240 0 0 $X=317210 $Y=46000
X1384 1 2 521 2 558 1 sky130_fd_sc_hd__clkbuf_4 $T=322000 40800 1 0 $X=321810 $Y=37840
X1385 1 2 521 2 559 1 sky130_fd_sc_hd__clkbuf_4 $T=322000 46240 1 0 $X=321810 $Y=43280
X1386 1 2 521 2 560 1 sky130_fd_sc_hd__clkbuf_4 $T=322000 51680 1 0 $X=321810 $Y=48720
X1387 1 2 521 2 561 1 sky130_fd_sc_hd__clkbuf_4 $T=322000 57120 1 0 $X=321810 $Y=54160
X1388 1 2 525 2 562 1 sky130_fd_sc_hd__clkbuf_4 $T=323840 35360 0 0 $X=323650 $Y=35120
X1389 1 2 525 2 563 1 sky130_fd_sc_hd__clkbuf_4 $T=323840 40800 0 0 $X=323650 $Y=40560
X1390 1 2 525 2 564 1 sky130_fd_sc_hd__clkbuf_4 $T=323840 51680 0 0 $X=323650 $Y=51440
X1391 1 2 525 2 565 1 sky130_fd_sc_hd__clkbuf_4 $T=323840 57120 0 0 $X=323650 $Y=56880
X1392 1 2 525 2 566 1 sky130_fd_sc_hd__clkbuf_4 $T=329820 46240 1 0 $X=329630 $Y=43280
X1393 1 2 525 2 567 1 sky130_fd_sc_hd__clkbuf_4 $T=330280 40800 0 0 $X=330090 $Y=40560
X1394 1 2 525 2 568 1 sky130_fd_sc_hd__clkbuf_4 $T=330280 51680 0 0 $X=330090 $Y=51440
X1395 1 2 525 2 569 1 sky130_fd_sc_hd__clkbuf_4 $T=333500 46240 0 0 $X=333310 $Y=46000
X1396 1 2 234 2 237 1 sky130_fd_sc_hd__clkbuf_16 $T=303140 35360 0 0 $X=302950 $Y=35120
X1397 1 2 235 2 504 1 sky130_fd_sc_hd__clkbuf_16 $T=306820 40800 1 0 $X=306630 $Y=37840
X1398 1 2 523 2 520 1 sky130_fd_sc_hd__clkbuf_16 $T=323380 46240 0 0 $X=323190 $Y=46000
X1399 1 2 395 149 129 2 440 1 sky130_fd_sc_hd__a21o_4 $T=176180 68000 0 0 $X=175990 $Y=67760
X1400 1 2 129 150 427 2 444 1 sky130_fd_sc_hd__a21o_4 $T=178020 78880 1 0 $X=177830 $Y=75920
X1401 1 2 395 145 148 2 441 1 sky130_fd_sc_hd__a21o_4 $T=178480 57120 1 0 $X=178290 $Y=54160
X1402 1 2 419 152 449 2 328 1 sky130_fd_sc_hd__a21o_4 $T=191820 62560 0 0 $X=191630 $Y=62320
X1403 1 2 456 137 198 2 479 1 sky130_fd_sc_hd__a21o_4 $T=251160 68000 1 0 $X=250970 $Y=65040
X1404 1 2 203 188 487 2 482 1 sky130_fd_sc_hd__a21o_4 $T=262660 51680 1 0 $X=262470 $Y=48720
X1405 1 2 203 188 492 2 491 1 sky130_fd_sc_hd__a21o_4 $T=270940 46240 0 0 $X=270750 $Y=46000
X1406 1 2 498 483 495 2 501 1 sky130_fd_sc_hd__a21o_4 $T=287500 57120 0 0 $X=287310 $Y=56880
X1407 1 2 498 483 510 2 511 1 sky130_fd_sc_hd__a21o_4 $T=301760 51680 0 0 $X=301570 $Y=51440
X1408 1 2 498 188 231 2 516 1 sky130_fd_sc_hd__a21o_4 $T=304980 73440 0 0 $X=304790 $Y=73200
X1409 1 2 498 188 514 2 517 1 sky130_fd_sc_hd__a21o_4 $T=305900 68000 1 0 $X=305710 $Y=65040
X1410 1 2 498 483 239 2 522 1 sky130_fd_sc_hd__a21o_4 $T=315560 68000 0 0 $X=315370 $Y=67760
X1411 1 2 8 10 ICV_39 $T=7820 46240 1 0 $X=7630 $Y=43280
X1412 1 2 7 8 ICV_39 $T=7820 51680 1 0 $X=7630 $Y=48720
X1413 1 2 7 8 ICV_39 $T=21160 46240 1 0 $X=20970 $Y=43280
X1414 1 2 349 355 ICV_39 $T=40020 62560 0 0 $X=39830 $Y=62320
X1415 1 2 329 38 ICV_39 $T=49220 51680 1 0 $X=49030 $Y=48720
X1416 1 2 67 382 ICV_39 $T=82800 35360 0 0 $X=82610 $Y=35120
X1417 1 2 64 384 ICV_39 $T=91080 40800 0 0 $X=90890 $Y=40560
X1418 1 2 51 396 ICV_39 $T=104880 40800 0 0 $X=104690 $Y=40560
X1419 1 2 96 406 ICV_39 $T=123280 51680 0 0 $X=123090 $Y=51440
X1420 1 2 430 411 ICV_39 $T=152260 68000 1 0 $X=152070 $Y=65040
X1421 1 2 112 133 ICV_39 $T=153180 78880 1 0 $X=152990 $Y=75920
X1422 1 2 136 431 ICV_39 $T=163300 68000 0 0 $X=163110 $Y=67760
X1423 1 2 436 429 ICV_39 $T=166980 57120 0 0 $X=166790 $Y=56880
X1424 1 2 410 385 ICV_39 $T=181700 46240 0 0 $X=181510 $Y=46000
X1425 1 2 449 152 ICV_39 $T=191820 62560 1 0 $X=191630 $Y=59600
X1426 1 2 170 120 ICV_39 $T=209300 78880 1 0 $X=209110 $Y=75920
X1427 1 2 194 470 ICV_39 $T=251160 68000 0 0 $X=250970 $Y=67760
X1428 1 2 202 474 ICV_39 $T=256220 73440 1 0 $X=256030 $Y=70480
X1429 1 2 8 519 ICV_39 $T=307280 57120 0 0 $X=307090 $Y=56880
X1430 1 2 142 444 145 419 435 2 442 1 sky130_fd_sc_hd__a32o_4 $T=175260 73440 0 0 $X=175070 $Y=73200
X1431 1 2 151 89 157 118 152 2 448 1 sky130_fd_sc_hd__a32o_4 $T=190900 78880 1 0 $X=190710 $Y=75920
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=36
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=10580 0 0 0 $X=10390 $Y=-240
X1 1 2 3 4 6 2 5 1 sky130_fd_sc_hd__dfrtp_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_42 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
** N=245 EP=199 IP=2688 FDC=4371
X0 1 2 Dpar a=554.335 p=693.97 m=1 $[nwdiode] $X=5330 $Y=10690 $D=191
X1 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=14905 $D=191
X2 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=20345 $D=191
X3 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=25785 $D=191
X4 1 2 Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=31225 $D=191
X5 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 13600 1 0 $X=5330 $Y=10640
X6 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 13600 0 0 $X=5330 $Y=13360
X7 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 19040 1 0 $X=5330 $Y=16080
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 19040 0 0 $X=5330 $Y=18800
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 24480 1 0 $X=5330 $Y=21520
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 24480 0 0 $X=5330 $Y=24240
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 29920 1 0 $X=5330 $Y=26960
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 29920 0 0 $X=5330 $Y=29680
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 35360 1 0 $X=5330 $Y=32400
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 35360 1 0 $X=6710 $Y=32400
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=22080 24480 0 0 $X=21890 $Y=24240
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 13600 0 0 $X=25570 $Y=13360
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 19040 1 0 $X=25570 $Y=16080
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=58420 13600 0 0 $X=58230 $Y=13360
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=58420 29920 0 0 $X=58230 $Y=29680
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=64860 35360 1 0 $X=64670 $Y=32400
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=82800 13600 0 0 $X=82610 $Y=13360
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=82800 29920 0 0 $X=82610 $Y=29680
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=87400 19040 1 0 $X=87210 $Y=16080
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=89700 13600 1 0 $X=89510 $Y=10640
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=104420 24480 1 0 $X=104230 $Y=21520
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=104420 29920 1 0 $X=104230 $Y=26960
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=112700 13600 0 0 $X=112510 $Y=13360
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 29920 1 0 $X=130450 $Y=26960
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=132480 24480 1 0 $X=132290 $Y=21520
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=140760 13600 0 0 $X=140570 $Y=13360
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 24480 0 0 $X=144250 $Y=24240
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=156400 35360 1 0 $X=156210 $Y=32400
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 35360 1 0 $X=158510 $Y=32400
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 24480 0 0 $X=174150 $Y=24240
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=175720 19040 1 0 $X=175530 $Y=16080
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=178020 19040 1 0 $X=177830 $Y=16080
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=195500 19040 0 0 $X=195310 $Y=18800
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=196880 29920 0 0 $X=196690 $Y=29680
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=197340 24480 1 0 $X=197150 $Y=21520
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=198720 13600 0 0 $X=198530 $Y=13360
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=209300 24480 1 0 $X=209110 $Y=21520
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=239660 13600 1 0 $X=239470 $Y=10640
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 24480 1 0 $X=242690 $Y=21520
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 29920 1 0 $X=242690 $Y=26960
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=253920 24480 1 0 $X=253730 $Y=21520
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=258520 13600 0 0 $X=258330 $Y=13360
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=258520 19040 0 0 $X=258330 $Y=18800
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286580 19040 0 0 $X=286390 $Y=18800
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=292100 24480 0 0 $X=291910 $Y=24240
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 29920 0 0 $X=314450 $Y=29680
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=318780 19040 1 0 $X=318590 $Y=16080
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 13600 0 180 $X=348950 $Y=10640
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 13600 1 180 $X=348950 $Y=13360
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 19040 0 180 $X=348950 $Y=16080
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 19040 1 180 $X=348950 $Y=18800
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 24480 0 180 $X=348950 $Y=21520
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 24480 1 180 $X=348950 $Y=24240
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 29920 0 180 $X=348950 $Y=26960
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 29920 1 180 $X=348950 $Y=29680
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350520 35360 0 180 $X=348950 $Y=32400
X113 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=23920 19040 0 0 $X=23730 $Y=18800
X114 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=25760 24480 1 0 $X=25570 $Y=21520
X115 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=35880 24480 0 0 $X=35690 $Y=24240
X116 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=39560 29920 1 0 $X=39370 $Y=26960
X117 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=43240 19040 1 0 $X=43050 $Y=16080
X118 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=48300 29920 1 0 $X=48110 $Y=26960
X119 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=48300 35360 1 0 $X=48110 $Y=32400
X120 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=65780 19040 0 0 $X=65590 $Y=18800
X121 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 13600 1 0 $X=72030 $Y=10640
X122 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=79120 13600 0 0 $X=78930 $Y=13360
X123 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=79120 29920 0 0 $X=78930 $Y=29680
X124 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100740 13600 1 0 $X=100550 $Y=10640
X125 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=109020 13600 0 0 $X=108830 $Y=13360
X126 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=123740 24480 0 0 $X=123550 $Y=24240
X127 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=126960 29920 1 0 $X=126770 $Y=26960
X128 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 35360 1 0 $X=128150 $Y=32400
X129 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=130180 29920 0 0 $X=129990 $Y=29680
X130 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 13600 1 0 $X=139650 $Y=10640
X131 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=155480 29920 1 0 $X=155290 $Y=26960
X132 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 19040 1 0 $X=156210 $Y=16080
X133 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 35360 1 0 $X=165410 $Y=32400
X134 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183540 29920 1 0 $X=183350 $Y=26960
X135 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=191820 19040 0 0 $X=191630 $Y=18800
X136 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=193660 24480 1 0 $X=193470 $Y=21520
X137 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194120 19040 1 0 $X=193930 $Y=16080
X138 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=202400 24480 0 0 $X=202210 $Y=24240
X139 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=207460 29920 0 0 $X=207270 $Y=29680
X140 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=207920 19040 0 0 $X=207730 $Y=18800
X141 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 13600 1 0 $X=210950 $Y=10640
X142 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211600 24480 1 0 $X=211410 $Y=21520
X143 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=224020 19040 1 0 $X=223830 $Y=16080
X144 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 24480 0 0 $X=230270 $Y=24240
X145 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 29920 0 0 $X=230270 $Y=29680
X146 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=235980 13600 0 0 $X=235790 $Y=13360
X147 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=239200 24480 1 0 $X=239010 $Y=21520
X148 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249780 35360 1 0 $X=249590 $Y=32400
X149 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=250240 24480 1 0 $X=250050 $Y=21520
X150 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=250700 19040 0 0 $X=250510 $Y=18800
X151 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=267720 24480 1 0 $X=267530 $Y=21520
X152 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=275540 13600 0 0 $X=275350 $Y=13360
X153 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278300 35360 1 0 $X=278110 $Y=32400
X154 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282440 24480 0 0 $X=282250 $Y=24240
X155 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=287040 13600 1 0 $X=286850 $Y=10640
X156 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 19040 1 0 $X=300650 $Y=16080
X157 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310040 29920 1 0 $X=309850 $Y=26960
X158 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 19040 0 0 $X=310310 $Y=18800
X159 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 29920 0 0 $X=310310 $Y=29680
X160 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 13600 0 0 $X=314450 $Y=13360
X161 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=316480 24480 1 0 $X=316290 $Y=21520
X162 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=320160 19040 0 0 $X=319970 $Y=18800
X163 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=323840 24480 1 0 $X=323650 $Y=21520
X164 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=330740 13600 0 0 $X=330550 $Y=13360
X165 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344540 19040 0 0 $X=344350 $Y=18800
X166 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345000 19040 1 0 $X=344810 $Y=16080
X167 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 13600 1 0 $X=12230 $Y=10640
X168 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=18400 19040 0 0 $X=18210 $Y=18800
X169 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=18400 29920 0 0 $X=18210 $Y=29680
X170 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=20240 13600 0 0 $X=20050 $Y=13360
X171 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=23920 29920 0 0 $X=23730 $Y=29680
X172 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25760 35360 1 0 $X=25570 $Y=32400
X173 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=34040 29920 1 0 $X=33850 $Y=26960
X174 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=37720 19040 1 0 $X=37530 $Y=16080
X175 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=37720 29920 0 0 $X=37530 $Y=29680
X176 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=45540 19040 0 0 $X=45350 $Y=18800
X177 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=47380 13600 0 0 $X=47190 $Y=13360
X178 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=53820 24480 1 0 $X=53630 $Y=21520
X179 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=53820 24480 0 0 $X=53630 $Y=24240
X180 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55200 29920 1 0 $X=55010 $Y=26960
X181 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=65780 24480 0 0 $X=65590 $Y=24240
X182 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=66240 19040 1 0 $X=66050 $Y=16080
X183 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=66700 13600 1 0 $X=66510 $Y=10640
X184 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=73600 13600 0 0 $X=73410 $Y=13360
X185 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81880 19040 1 0 $X=81690 $Y=16080
X186 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81880 29920 1 0 $X=81690 $Y=26960
X187 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=82800 13600 1 0 $X=82610 $Y=10640
X188 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=88320 35360 1 0 $X=88130 $Y=32400
X189 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=95220 13600 1 0 $X=95030 $Y=10640
X190 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=95220 24480 1 0 $X=95030 $Y=21520
X191 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97980 35360 1 0 $X=97790 $Y=32400
X192 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=102580 29920 0 0 $X=102390 $Y=29680
X193 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=103040 19040 0 0 $X=102850 $Y=18800
X194 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=108560 19040 0 0 $X=108370 $Y=18800
X195 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=111780 24480 0 0 $X=111590 $Y=24240
X196 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=124660 19040 1 0 $X=124470 $Y=16080
X197 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=129720 13600 0 0 $X=129530 $Y=13360
X198 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=135240 13600 0 0 $X=135050 $Y=13360
X199 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=138000 19040 1 0 $X=137810 $Y=16080
X200 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=138000 35360 1 0 $X=137810 $Y=32400
X201 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=149960 29920 1 0 $X=149770 $Y=26960
X202 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=151800 24480 0 0 $X=151610 $Y=24240
X203 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=155940 13600 1 0 $X=155750 $Y=10640
X204 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=157320 24480 0 0 $X=157130 $Y=24240
X205 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=162840 24480 0 0 $X=162650 $Y=24240
X206 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=166060 29920 1 0 $X=165870 $Y=26960
X207 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=168360 24480 0 0 $X=168170 $Y=24240
X208 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=171580 29920 1 0 $X=171390 $Y=26960
X209 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=179860 35360 1 0 $X=179670 $Y=32400
X210 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=184460 13600 1 0 $X=184270 $Y=10640
X211 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=187680 13600 0 0 $X=187490 $Y=13360
X212 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=193200 13600 0 0 $X=193010 $Y=13360
X213 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=206080 13600 0 0 $X=205890 $Y=13360
X214 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210680 35360 1 0 $X=210490 $Y=32400
X215 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=220340 24480 1 0 $X=220150 $Y=21520
X216 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=245180 19040 0 0 $X=244990 $Y=18800
X217 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=264040 29920 0 0 $X=263850 $Y=29680
X218 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=269560 29920 0 0 $X=269370 $Y=29680
X219 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=275080 29920 0 0 $X=274890 $Y=29680
X220 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=285660 29920 1 0 $X=285470 $Y=26960
X221 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=290720 24480 1 0 $X=290530 $Y=21520
X222 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=291180 29920 1 0 $X=290990 $Y=26960
X223 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=304520 29920 1 0 $X=304330 $Y=26960
X224 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=312800 13600 1 0 $X=312610 $Y=10640
X225 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=327060 13600 1 0 $X=326870 $Y=10640
X226 1 2 ICV_2 $T=19780 13600 1 0 $X=19590 $Y=10640
X227 1 2 ICV_2 $T=19780 19040 1 0 $X=19590 $Y=16080
X228 1 2 ICV_2 $T=19780 24480 1 0 $X=19590 $Y=21520
X229 1 2 ICV_2 $T=19780 35360 1 0 $X=19590 $Y=32400
X230 1 2 ICV_2 $T=47840 19040 1 0 $X=47650 $Y=16080
X231 1 2 ICV_2 $T=47840 24480 1 0 $X=47650 $Y=21520
X232 1 2 ICV_2 $T=48300 13600 1 0 $X=48110 $Y=10640
X233 1 2 ICV_2 $T=75900 29920 1 0 $X=75710 $Y=26960
X234 1 2 ICV_2 $T=76820 13600 1 0 $X=76630 $Y=10640
X235 1 2 ICV_2 $T=103960 35360 1 0 $X=103770 $Y=32400
X236 1 2 ICV_2 $T=105340 13600 1 0 $X=105150 $Y=10640
X237 1 2 ICV_2 $T=117760 24480 0 0 $X=117570 $Y=24240
X238 1 2 ICV_2 $T=119600 13600 1 0 $X=119410 $Y=10640
X239 1 2 ICV_2 $T=132020 19040 1 0 $X=131830 $Y=16080
X240 1 2 ICV_2 $T=132020 35360 1 0 $X=131830 $Y=32400
X241 1 2 ICV_2 $T=133860 13600 1 0 $X=133670 $Y=10640
X242 1 2 ICV_2 $T=145820 24480 0 0 $X=145630 $Y=24240
X243 1 2 ICV_2 $T=160080 24480 1 0 $X=159890 $Y=21520
X244 1 2 ICV_2 $T=160080 29920 1 0 $X=159890 $Y=26960
X245 1 2 ICV_2 $T=162380 13600 1 0 $X=162190 $Y=10640
X246 1 2 ICV_2 $T=173880 29920 0 0 $X=173690 $Y=29680
X247 1 2 ICV_2 $T=188140 19040 1 0 $X=187950 $Y=16080
X248 1 2 ICV_2 $T=190900 13600 1 0 $X=190710 $Y=10640
X249 1 2 ICV_2 $T=201940 19040 0 0 $X=201750 $Y=18800
X250 1 2 ICV_2 $T=205160 13600 1 0 $X=204970 $Y=10640
X251 1 2 ICV_2 $T=219420 13600 1 0 $X=219230 $Y=10640
X252 1 2 ICV_2 $T=233680 13600 1 0 $X=233490 $Y=10640
X253 1 2 ICV_2 $T=244260 24480 1 0 $X=244070 $Y=21520
X254 1 2 ICV_2 $T=244260 29920 1 0 $X=244070 $Y=26960
X255 1 2 ICV_2 $T=247940 13600 1 0 $X=247750 $Y=10640
X256 1 2 ICV_2 $T=258060 29920 0 0 $X=257870 $Y=29680
X257 1 2 ICV_2 $T=272320 19040 1 0 $X=272130 $Y=16080
X258 1 2 ICV_2 $T=272320 35360 1 0 $X=272130 $Y=32400
X259 1 2 ICV_2 $T=286120 13600 0 0 $X=285930 $Y=13360
X260 1 2 ICV_2 $T=286120 24480 0 0 $X=285930 $Y=24240
X261 1 2 ICV_2 $T=286120 29920 0 0 $X=285930 $Y=29680
X262 1 2 ICV_2 $T=290720 13600 1 0 $X=290530 $Y=10640
X263 1 2 ICV_2 $T=314180 19040 0 0 $X=313990 $Y=18800
X264 1 2 ICV_2 $T=328440 35360 1 0 $X=328250 $Y=32400
X265 1 2 ICV_2 $T=333500 13600 1 0 $X=333310 $Y=10640
X266 1 2 ICV_2 $T=342240 13600 0 0 $X=342050 $Y=13360
X267 1 2 ICV_2 $T=342240 24480 0 0 $X=342050 $Y=24240
X268 1 2 ICV_2 $T=342240 29920 0 0 $X=342050 $Y=29680
X269 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 13600 1 0 $X=17750 $Y=10640
X270 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 19040 1 0 $X=17750 $Y=16080
X271 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 24480 1 0 $X=17750 $Y=21520
X272 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 29920 1 0 $X=17750 $Y=26960
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=29440 29920 0 0 $X=29250 $Y=29680
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31280 35360 1 0 $X=31090 $Y=32400
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34500 13600 1 0 $X=34310 $Y=10640
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=44160 35360 1 0 $X=43970 $Y=32400
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=53820 19040 1 0 $X=53630 $Y=16080
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59340 24480 1 0 $X=59150 $Y=21520
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 29920 0 0 $X=61910 $Y=29680
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=74520 29920 0 0 $X=74330 $Y=29680
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=86020 24480 0 0 $X=85830 $Y=24240
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=90160 19040 0 0 $X=89970 $Y=18800
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=97520 24480 0 0 $X=97330 $Y=24240
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=114080 29920 0 0 $X=113890 $Y=29680
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 19040 1 0 $X=115730 $Y=16080
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 19040 0 0 $X=118030 $Y=18800
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=123740 29920 1 0 $X=123550 $Y=26960
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=130180 19040 1 0 $X=129990 $Y=16080
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=140300 29920 0 0 $X=140110 $Y=29680
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 35360 1 0 $X=143330 $Y=32400
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=166060 24480 1 0 $X=165870 $Y=21520
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=166980 29920 0 0 $X=166790 $Y=29680
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 29920 0 0 $X=171850 $Y=29680
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=177100 29920 1 0 $X=176910 $Y=26960
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=185840 19040 1 0 $X=185650 $Y=16080
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 24480 1 0 $X=186110 $Y=21520
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=199640 19040 0 0 $X=199450 $Y=18800
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=212520 29920 1 0 $X=212330 $Y=26960
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226320 13600 0 0 $X=226130 $Y=13360
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226320 19040 0 0 $X=226130 $Y=18800
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230460 19040 0 0 $X=230270 $Y=18800
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=240580 19040 1 0 $X=240390 $Y=16080
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=262660 13600 1 0 $X=262470 $Y=10640
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=262660 19040 1 0 $X=262470 $Y=16080
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=272780 29920 1 0 $X=272590 $Y=26960
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=292100 29920 0 0 $X=291910 $Y=29680
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=303140 13600 1 0 $X=302950 $Y=10640
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 35360 1 0 $X=325950 $Y=32400
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 19040 1 0 $X=326410 $Y=16080
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=332580 24480 1 0 $X=332390 $Y=21520
X311 1 19 sky130_fd_sc_hd__diode_2 $T=34960 24480 0 0 $X=34770 $Y=24240
X312 1 7 sky130_fd_sc_hd__diode_2 $T=57500 13600 0 0 $X=57310 $Y=13360
X313 1 29 sky130_fd_sc_hd__diode_2 $T=57500 29920 0 0 $X=57310 $Y=29680
X314 1 7 sky130_fd_sc_hd__diode_2 $T=63940 35360 1 0 $X=63750 $Y=32400
X315 1 7 sky130_fd_sc_hd__diode_2 $T=72220 19040 1 0 $X=72030 $Y=16080
X316 1 46 sky130_fd_sc_hd__diode_2 $T=83720 19040 0 0 $X=83530 $Y=18800
X317 1 7 sky130_fd_sc_hd__diode_2 $T=88780 13600 1 0 $X=88590 $Y=10640
X318 1 61 sky130_fd_sc_hd__diode_2 $T=108100 13600 0 0 $X=107910 $Y=13360
X319 1 44 sky130_fd_sc_hd__diode_2 $T=108100 29920 0 0 $X=107910 $Y=29680
X320 1 7 sky130_fd_sc_hd__diode_2 $T=118220 19040 1 0 $X=118030 $Y=16080
X321 1 70 sky130_fd_sc_hd__diode_2 $T=118680 35360 1 0 $X=118490 $Y=32400
X322 1 73 sky130_fd_sc_hd__diode_2 $T=124200 29920 0 0 $X=124010 $Y=29680
X323 1 74 sky130_fd_sc_hd__diode_2 $T=126040 29920 1 0 $X=125850 $Y=26960
X324 1 75 sky130_fd_sc_hd__diode_2 $T=127420 35360 1 0 $X=127230 $Y=32400
X325 1 79 sky130_fd_sc_hd__diode_2 $T=134320 29920 0 0 $X=134130 $Y=29680
X326 1 93 sky130_fd_sc_hd__diode_2 $T=157780 35360 1 0 $X=157590 $Y=32400
X327 1 7 sky130_fd_sc_hd__diode_2 $T=177100 19040 1 0 $X=176910 $Y=16080
X328 1 225 sky130_fd_sc_hd__diode_2 $T=182620 29920 1 0 $X=182430 $Y=26960
X329 1 224 sky130_fd_sc_hd__diode_2 $T=190900 19040 0 0 $X=190710 $Y=18800
X330 1 112 sky130_fd_sc_hd__diode_2 $T=201020 35360 1 0 $X=200830 $Y=32400
X331 1 226 sky130_fd_sc_hd__diode_2 $T=210680 24480 1 0 $X=210490 $Y=21520
X332 1 7 sky130_fd_sc_hd__diode_2 $T=215740 13600 1 0 $X=215550 $Y=10640
X333 1 132 sky130_fd_sc_hd__diode_2 $T=235060 13600 0 0 $X=234870 $Y=13360
X334 1 151 sky130_fd_sc_hd__diode_2 $T=268180 35360 1 0 $X=267990 $Y=32400
X335 1 7 sky130_fd_sc_hd__diode_2 $T=270940 24480 0 0 $X=270750 $Y=24240
X336 1 159 sky130_fd_sc_hd__diode_2 $T=281520 24480 0 0 $X=281330 $Y=24240
X337 1 7 sky130_fd_sc_hd__diode_2 $T=284280 29920 0 0 $X=284090 $Y=29680
X338 1 170 sky130_fd_sc_hd__diode_2 $T=296700 19040 1 0 $X=296510 $Y=16080
X339 1 177 sky130_fd_sc_hd__diode_2 $T=309580 19040 0 0 $X=309390 $Y=18800
X340 1 194 sky130_fd_sc_hd__diode_2 $T=338100 13600 0 0 $X=337910 $Y=13360
X341 1 195 sky130_fd_sc_hd__diode_2 $T=338100 29920 0 0 $X=337910 $Y=29680
X342 1 7 sky130_fd_sc_hd__diode_2 $T=343620 19040 0 0 $X=343430 $Y=18800
X343 1 2 15 ICV_4 $T=30820 13600 0 0 $X=30630 $Y=13360
X344 1 2 7 ICV_4 $T=43240 29920 1 0 $X=43050 $Y=26960
X345 1 2 42 ICV_4 $T=73140 24480 1 0 $X=72950 $Y=21520
X346 1 2 7 ICV_4 $T=101200 24480 1 0 $X=101010 $Y=21520
X347 1 2 59 ICV_4 $T=101200 29920 1 0 $X=101010 $Y=26960
X348 1 2 7 ICV_4 $T=179400 29920 1 0 $X=179210 $Y=26960
X349 1 2 112 ICV_4 $T=194580 35360 1 0 $X=194390 $Y=32400
X350 1 2 115 ICV_4 $T=198720 19040 1 0 $X=198530 $Y=16080
X351 1 2 3 ICV_4 $T=244720 13600 1 0 $X=244530 $Y=10640
X352 1 2 7 ICV_4 $T=253000 24480 0 0 $X=252810 $Y=24240
X353 1 2 7 ICV_4 $T=257140 19040 1 0 $X=256950 $Y=16080
X354 1 2 147 ICV_4 $T=259900 13600 0 0 $X=259710 $Y=13360
X355 1 2 7 ICV_4 $T=283360 13600 0 0 $X=283170 $Y=13360
X356 1 2 7 ICV_4 $T=297160 24480 1 0 $X=296970 $Y=21520
X357 1 2 189 ICV_4 $T=329820 19040 1 0 $X=329630 $Y=16080
X358 1 2 3 ICV_4 $T=339480 19040 0 0 $X=339290 $Y=18800
X359 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 13600 1 0 $X=6710 $Y=10640
X360 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=20240 29920 1 0 $X=20050 $Y=26960
X361 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 35360 1 0 $X=72490 $Y=32400
X362 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 19040 1 0 $X=72950 $Y=16080
X363 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=76360 19040 1 0 $X=76170 $Y=16080
X364 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=76360 24480 1 0 $X=76170 $Y=21520
X365 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=81420 35360 1 0 $X=81230 $Y=32400
X366 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=84640 19040 0 0 $X=84450 $Y=18800
X367 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=89700 24480 1 0 $X=89510 $Y=21520
X368 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=98440 29920 1 0 $X=98250 $Y=26960
X369 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101660 13600 0 0 $X=101470 $Y=13360
X370 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=119140 19040 1 0 $X=118950 $Y=16080
X371 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=119600 35360 1 0 $X=119410 $Y=32400
X372 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=127420 24480 1 0 $X=127230 $Y=21520
X373 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 19040 0 0 $X=132290 $Y=18800
X374 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 29920 1 0 $X=132290 $Y=26960
X375 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 24480 1 0 $X=146090 $Y=21520
X376 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157780 13600 0 0 $X=157590 $Y=13360
X377 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157780 29920 0 0 $X=157590 $Y=29680
X378 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=170660 13600 0 0 $X=170470 $Y=13360
X379 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=174340 19040 0 0 $X=174150 $Y=18800
X380 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=200100 29920 1 0 $X=199910 $Y=26960
X381 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=205620 29920 1 0 $X=205430 $Y=26960
X382 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 13600 1 0 $X=216470 $Y=10640
X383 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=264960 35360 1 0 $X=264770 $Y=32400
X384 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269100 29920 1 0 $X=268910 $Y=26960
X385 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269100 35360 1 0 $X=268910 $Y=32400
X386 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=270480 19040 0 0 $X=270290 $Y=18800
X387 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=271400 13600 1 0 $X=271210 $Y=10640
X388 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=278300 19040 1 0 $X=278110 $Y=16080
X389 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=292100 13600 0 0 $X=291910 $Y=13360
X390 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297620 19040 1 0 $X=297430 $Y=16080
X391 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=310960 13600 0 0 $X=310770 $Y=13360
X392 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339020 13600 0 0 $X=338830 $Y=13360
X393 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339020 24480 0 0 $X=338830 $Y=24240
X394 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339020 29920 0 0 $X=338830 $Y=29680
X395 1 3 7 ICV_7 $T=7820 19040 1 0 $X=7630 $Y=16080
X396 1 3 7 ICV_7 $T=7820 24480 1 0 $X=7630 $Y=21520
X397 1 3 7 ICV_7 $T=7820 29920 1 0 $X=7630 $Y=26960
X398 1 3 8 ICV_7 $T=8280 35360 1 0 $X=8090 $Y=32400
X399 1 7 9 ICV_7 $T=9660 13600 1 0 $X=9470 $Y=10640
X400 1 3 7 ICV_7 $T=23460 24480 0 0 $X=23270 $Y=24240
X401 1 3 7 ICV_7 $T=27140 13600 0 0 $X=26950 $Y=13360
X402 1 7 3 ICV_7 $T=28060 19040 0 0 $X=27870 $Y=18800
X403 1 16 7 ICV_7 $T=29900 24480 1 0 $X=29710 $Y=21520
X404 1 3 7 ICV_7 $T=34960 29920 0 0 $X=34770 $Y=29680
X405 1 7 21 ICV_7 $T=36800 13600 1 0 $X=36610 $Y=10640
X406 1 22 3 ICV_7 $T=39560 24480 0 0 $X=39370 $Y=24240
X407 1 3 7 ICV_7 $T=52440 29920 1 0 $X=52250 $Y=26960
X408 1 30 3 ICV_7 $T=53820 13600 0 0 $X=53630 $Y=13360
X409 1 3 7 ICV_7 $T=63020 19040 0 0 $X=62830 $Y=18800
X410 1 3 7 ICV_7 $T=63020 24480 0 0 $X=62830 $Y=24240
X411 1 7 36 ICV_7 $T=63940 13600 1 0 $X=63750 $Y=10640
X412 1 220 7 ICV_7 $T=71760 24480 0 0 $X=71570 $Y=24240
X413 1 44 45 ICV_7 $T=76360 29920 0 0 $X=76170 $Y=29680
X414 1 3 7 ICV_7 $T=79120 19040 1 0 $X=78930 $Y=16080
X415 1 48 3 ICV_7 $T=84180 13600 0 0 $X=83990 $Y=13360
X416 1 44 50 ICV_7 $T=84180 29920 0 0 $X=83990 $Y=29680
X417 1 7 54 ICV_7 $T=92460 13600 1 0 $X=92270 $Y=10640
X418 1 3 7 ICV_7 $T=92460 24480 1 0 $X=92270 $Y=21520
X419 1 3 7 ICV_7 $T=104420 13600 0 0 $X=104230 $Y=13360
X420 1 7 62 ICV_7 $T=105800 24480 1 0 $X=105610 $Y=21520
X421 1 63 65 ICV_7 $T=109940 35360 1 0 $X=109750 $Y=32400
X422 1 66 3 ICV_7 $T=114080 13600 0 0 $X=113890 $Y=13360
X423 1 222 7 ICV_7 $T=114080 19040 0 0 $X=113890 $Y=18800
X424 1 7 72 ICV_7 $T=121900 19040 1 0 $X=121710 $Y=16080
X425 1 3 7 ICV_7 $T=135700 19040 0 0 $X=135510 $Y=18800
X426 1 3 7 ICV_7 $T=141680 24480 0 0 $X=141490 $Y=24240
X427 1 7 3 ICV_7 $T=142140 13600 0 0 $X=141950 $Y=13360
X428 1 82 7 ICV_7 $T=142140 29920 0 0 $X=141950 $Y=29680
X429 1 83 3 ICV_7 $T=144440 13600 1 0 $X=144250 $Y=10640
X430 1 7 87 ICV_7 $T=147200 29920 1 0 $X=147010 $Y=26960
X431 1 7 88 ICV_7 $T=149040 24480 1 0 $X=148850 $Y=21520
X432 1 3 7 ICV_7 $T=160540 13600 0 0 $X=160350 $Y=13360
X433 1 3 7 ICV_7 $T=168360 19040 0 0 $X=168170 $Y=18800
X434 1 7 98 ICV_7 $T=169280 29920 0 0 $X=169090 $Y=29680
X435 1 224 3 ICV_7 $T=175720 24480 0 0 $X=175530 $Y=24240
X436 1 3 7 ICV_7 $T=190900 24480 0 0 $X=190710 $Y=24240
X437 1 109 110 ICV_7 $T=194120 29920 0 0 $X=193930 $Y=29680
X438 1 7 3 ICV_7 $T=196880 19040 0 0 $X=196690 $Y=18800
X439 1 113 104 ICV_7 $T=197340 35360 1 0 $X=197150 $Y=32400
X440 1 114 109 ICV_7 $T=198260 29920 0 0 $X=198070 $Y=29680
X441 1 109 118 ICV_7 $T=202860 29920 1 0 $X=202670 $Y=26960
X442 1 3 7 ICV_7 $T=203320 13600 0 0 $X=203130 $Y=13360
X443 1 228 7 ICV_7 $T=207000 24480 0 0 $X=206810 $Y=24240
X444 1 119 121 ICV_7 $T=207920 35360 1 0 $X=207730 $Y=32400
X445 1 122 3 ICV_7 $T=212060 13600 0 0 $X=211870 $Y=13360
X446 1 7 3 ICV_7 $T=212060 19040 0 0 $X=211870 $Y=18800
X447 1 124 7 ICV_7 $T=212060 29920 0 0 $X=211870 $Y=29680
X448 1 7 227 ICV_7 $T=217580 24480 1 0 $X=217390 $Y=21520
X449 1 3 7 ICV_7 $T=231380 13600 0 0 $X=231190 $Y=13360
X450 1 7 3 ICV_7 $T=240120 13600 0 0 $X=239930 $Y=13360
X451 1 137 7 ICV_7 $T=241040 13600 1 0 $X=240850 $Y=10640
X452 1 229 3 ICV_7 $T=249320 24480 0 0 $X=249130 $Y=24240
X453 1 143 3 ICV_7 $T=254380 19040 0 0 $X=254190 $Y=18800
X454 1 7 146 ICV_7 $T=254380 29920 0 0 $X=254190 $Y=29680
X455 1 3 7 ICV_7 $T=259900 19040 1 0 $X=259710 $Y=16080
X456 1 3 7 ICV_7 $T=273700 19040 0 0 $X=273510 $Y=18800
X457 1 3 158 ICV_7 $T=277840 24480 0 0 $X=277650 $Y=24240
X458 1 160 3 ICV_7 $T=279680 13600 0 0 $X=279490 $Y=13360
X459 1 161 3 ICV_7 $T=280600 29920 0 0 $X=280410 $Y=29680
X460 1 3 165 ICV_7 $T=287960 24480 1 0 $X=287770 $Y=21520
X461 1 168 3 ICV_7 $T=293480 24480 0 0 $X=293290 $Y=24240
X462 1 169 3 ICV_7 $T=294400 29920 0 0 $X=294210 $Y=29680
X463 1 171 7 ICV_7 $T=296700 29920 1 0 $X=296510 $Y=26960
X464 1 164 7 ICV_7 $T=296700 35360 1 0 $X=296510 $Y=32400
X465 1 3 7 ICV_7 $T=305900 19040 0 0 $X=305710 $Y=18800
X466 1 3 175 ICV_7 $T=308200 13600 0 0 $X=308010 $Y=13360
X467 1 3 7 ICV_7 $T=315560 24480 0 0 $X=315370 $Y=24240
X468 1 185 3 ICV_7 $T=316020 29920 0 0 $X=315830 $Y=29680
X469 1 7 187 ICV_7 $T=321080 24480 1 0 $X=320890 $Y=21520
X470 1 7 3 ICV_7 $T=324300 19040 0 0 $X=324110 $Y=18800
X471 1 7 228 ICV_7 $T=329820 24480 1 0 $X=329630 $Y=21520
X472 1 3 7 ICV_7 $T=334420 13600 0 0 $X=334230 $Y=13360
X473 1 3 7 ICV_7 $T=334420 29920 0 0 $X=334230 $Y=29680
X474 1 2 3 4 7 2 10 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 19040 0 0 $X=7630 $Y=18800
X475 1 2 3 6 7 2 12 1 sky130_fd_sc_hd__dfrtp_4 $T=7820 29920 0 0 $X=7630 $Y=29680
X476 1 2 3 14 7 2 18 1 sky130_fd_sc_hd__dfrtp_4 $T=23460 29920 1 0 $X=23270 $Y=26960
X477 1 2 3 15 7 2 20 1 sky130_fd_sc_hd__dfrtp_4 $T=27140 19040 1 0 $X=26950 $Y=16080
X478 1 2 3 17 7 2 24 1 sky130_fd_sc_hd__dfrtp_4 $T=33580 35360 1 0 $X=33390 $Y=32400
X479 1 2 3 19 7 2 25 1 sky130_fd_sc_hd__dfrtp_4 $T=34960 19040 0 0 $X=34770 $Y=18800
X480 1 2 3 22 7 2 28 1 sky130_fd_sc_hd__dfrtp_4 $T=43240 24480 0 0 $X=43050 $Y=24240
X481 1 2 3 29 7 2 35 1 sky130_fd_sc_hd__dfrtp_4 $T=52440 35360 1 0 $X=52250 $Y=32400
X482 1 2 3 30 7 2 37 1 sky130_fd_sc_hd__dfrtp_4 $T=55660 19040 1 0 $X=55470 $Y=16080
X483 1 2 3 32 7 2 39 1 sky130_fd_sc_hd__dfrtp_4 $T=61640 24480 1 0 $X=61450 $Y=21520
X484 1 2 3 36 7 2 41 1 sky130_fd_sc_hd__dfrtp_4 $T=63020 13600 0 0 $X=62830 $Y=13360
X485 1 2 231 34 7 2 43 1 sky130_fd_sc_hd__dfrtp_4 $T=63940 29920 0 0 $X=63750 $Y=29680
X486 1 2 232 220 7 2 49 1 sky130_fd_sc_hd__dfrtp_4 $T=75440 24480 0 0 $X=75250 $Y=24240
X487 1 2 3 46 7 2 52 1 sky130_fd_sc_hd__dfrtp_4 $T=79120 24480 1 0 $X=78930 $Y=21520
X488 1 2 233 221 7 2 56 1 sky130_fd_sc_hd__dfrtp_4 $T=87860 29920 1 0 $X=87670 $Y=26960
X489 1 2 3 54 7 2 58 1 sky130_fd_sc_hd__dfrtp_4 $T=91080 13600 0 0 $X=90890 $Y=13360
X490 1 2 3 51 7 2 60 1 sky130_fd_sc_hd__dfrtp_4 $T=92460 19040 0 0 $X=92270 $Y=18800
X491 1 2 3 61 7 2 67 1 sky130_fd_sc_hd__dfrtp_4 $T=105340 19040 1 0 $X=105150 $Y=16080
X492 1 2 234 62 7 2 68 1 sky130_fd_sc_hd__dfrtp_4 $T=105800 29920 1 0 $X=105610 $Y=26960
X493 1 2 235 222 7 2 73 1 sky130_fd_sc_hd__dfrtp_4 $T=116840 24480 1 0 $X=116650 $Y=21520
X494 1 2 3 66 7 2 76 1 sky130_fd_sc_hd__dfrtp_4 $T=119140 13600 0 0 $X=118950 $Y=13360
X495 1 2 3 78 7 2 86 1 sky130_fd_sc_hd__dfrtp_4 $T=135700 29920 1 0 $X=135510 $Y=26960
X496 1 2 236 82 7 2 90 1 sky130_fd_sc_hd__dfrtp_4 $T=145820 35360 1 0 $X=145630 $Y=32400
X497 1 2 3 83 7 2 91 1 sky130_fd_sc_hd__dfrtp_4 $T=147200 13600 0 0 $X=147010 $Y=13360
X498 1 2 237 87 7 2 92 1 sky130_fd_sc_hd__dfrtp_4 $T=147200 29920 0 0 $X=147010 $Y=29680
X499 1 2 3 97 7 2 101 1 sky130_fd_sc_hd__dfrtp_4 $T=168360 24480 1 0 $X=168170 $Y=21520
X500 1 2 238 98 7 2 102 1 sky130_fd_sc_hd__dfrtp_4 $T=169280 35360 1 0 $X=169090 $Y=32400
X501 1 2 3 224 7 2 107 1 sky130_fd_sc_hd__dfrtp_4 $T=179400 24480 0 0 $X=179210 $Y=24240
X502 1 2 3 108 7 2 116 1 sky130_fd_sc_hd__dfrtp_4 $T=189520 29920 1 0 $X=189330 $Y=26960
X503 1 2 3 115 7 2 120 1 sky130_fd_sc_hd__dfrtp_4 $T=198720 24480 1 0 $X=198530 $Y=21520
X504 1 2 239 226 7 2 125 1 sky130_fd_sc_hd__dfrtp_4 $T=210680 24480 0 0 $X=210490 $Y=24240
X505 1 2 3 122 7 2 128 1 sky130_fd_sc_hd__dfrtp_4 $T=215740 13600 0 0 $X=215550 $Y=13360
X506 1 2 3 126 7 2 129 1 sky130_fd_sc_hd__dfrtp_4 $T=215740 19040 0 0 $X=215550 $Y=18800
X507 1 2 240 227 7 2 228 1 sky130_fd_sc_hd__dfrtp_4 $T=217580 29920 1 0 $X=217390 $Y=26960
X508 1 2 3 137 7 2 144 1 sky130_fd_sc_hd__dfrtp_4 $T=245640 19040 1 0 $X=245450 $Y=16080
X509 1 2 3 229 7 2 148 1 sky130_fd_sc_hd__dfrtp_4 $T=251160 29920 1 0 $X=250970 $Y=26960
X510 1 2 241 146 7 2 33 1 sky130_fd_sc_hd__dfrtp_4 $T=254380 35360 1 0 $X=254190 $Y=32400
X511 1 2 3 145 7 2 152 1 sky130_fd_sc_hd__dfrtp_4 $T=259440 24480 0 0 $X=259250 $Y=24240
X512 1 2 3 147 7 2 153 1 sky130_fd_sc_hd__dfrtp_4 $T=259900 19040 0 0 $X=259710 $Y=18800
X513 1 2 3 159 7 2 163 1 sky130_fd_sc_hd__dfrtp_4 $T=275080 29920 1 0 $X=274890 $Y=26960
X514 1 2 3 165 7 2 172 1 sky130_fd_sc_hd__dfrtp_4 $T=287960 19040 0 0 $X=287770 $Y=18800
X515 1 2 3 171 7 2 180 1 sky130_fd_sc_hd__dfrtp_4 $T=301760 35360 1 0 $X=301570 $Y=32400
X516 1 2 3 189 7 2 196 1 sky130_fd_sc_hd__dfrtp_4 $T=327980 19040 0 0 $X=327790 $Y=18800
X517 1 2 3 228 7 2 197 1 sky130_fd_sc_hd__dfrtp_4 $T=329820 29920 1 0 $X=329630 $Y=26960
X518 1 2 ICV_9 $T=11040 35360 1 0 $X=10850 $Y=32400
X519 1 2 ICV_9 $T=25760 13600 1 0 $X=25570 $Y=10640
X520 1 2 ICV_9 $T=39560 13600 1 0 $X=39370 $Y=10640
X521 1 2 ICV_9 $T=51060 19040 0 0 $X=50870 $Y=18800
X522 1 2 ICV_9 $T=54280 13600 1 0 $X=54090 $Y=10640
X523 1 2 ICV_9 $T=108560 24480 1 0 $X=108370 $Y=21520
X524 1 2 ICV_9 $T=111320 13600 1 0 $X=111130 $Y=10640
X525 1 2 ICV_9 $T=125580 13600 1 0 $X=125390 $Y=10640
X526 1 2 ICV_9 $T=151800 24480 1 0 $X=151610 $Y=21520
X527 1 2 ICV_9 $T=159620 19040 0 0 $X=159430 $Y=18800
X528 1 2 ICV_9 $T=168360 13600 1 0 $X=168170 $Y=10640
X529 1 2 ICV_9 $T=196880 13600 1 0 $X=196690 $Y=10640
X530 1 2 ICV_9 $T=221260 24480 0 0 $X=221070 $Y=24240
X531 1 2 ICV_9 $T=225400 13600 1 0 $X=225210 $Y=10640
X532 1 2 ICV_9 $T=228160 29920 1 0 $X=227970 $Y=26960
X533 1 2 ICV_9 $T=229080 35360 1 0 $X=228890 $Y=32400
X534 1 2 ICV_9 $T=241040 24480 0 0 $X=240850 $Y=24240
X535 1 2 ICV_9 $T=253920 13600 1 0 $X=253730 $Y=10640
X536 1 2 ICV_9 $T=339480 13600 1 0 $X=339290 $Y=10640
X537 1 2 ICV_9 $T=340400 29920 1 0 $X=340210 $Y=26960
X538 1 3 ICV_15 $T=31740 19040 0 0 $X=31550 $Y=18800
X539 1 17 ICV_15 $T=31740 29920 0 0 $X=31550 $Y=29680
X540 1 7 ICV_15 $T=46000 29920 1 0 $X=45810 $Y=26960
X541 1 26 ICV_15 $T=46000 35360 1 0 $X=45810 $Y=32400
X542 1 3 ICV_15 $T=59800 13600 0 0 $X=59610 $Y=13360
X543 1 32 ICV_15 $T=59800 19040 0 0 $X=59610 $Y=18800
X544 1 33 ICV_15 $T=59800 24480 0 0 $X=59610 $Y=24240
X545 1 34 ICV_15 $T=59800 29920 0 0 $X=59610 $Y=29680
X546 1 3 ICV_15 $T=87860 13600 0 0 $X=87670 $Y=13360
X547 1 51 ICV_15 $T=87860 19040 0 0 $X=87670 $Y=18800
X548 1 7 ICV_15 $T=87860 24480 0 0 $X=87670 $Y=24240
X549 1 49 ICV_15 $T=87860 29920 0 0 $X=87670 $Y=29680
X550 1 68 ICV_15 $T=115920 29920 0 0 $X=115730 $Y=29680
X551 1 223 ICV_15 $T=130180 24480 1 0 $X=129990 $Y=21520
X552 1 97 ICV_15 $T=172040 19040 0 0 $X=171850 $Y=18800
X553 1 104 ICV_15 $T=186300 35360 1 0 $X=186110 $Y=32400
X554 1 117 ICV_15 $T=200100 13600 0 0 $X=199910 $Y=13360
X555 1 125 ICV_15 $T=214360 29920 1 0 $X=214170 $Y=26960
X556 1 131 ICV_15 $T=228160 13600 0 0 $X=227970 $Y=13360
X557 1 3 ICV_15 $T=228160 19040 0 0 $X=227970 $Y=18800
X558 1 138 ICV_15 $T=242420 19040 1 0 $X=242230 $Y=16080
X559 1 3 ICV_15 $T=256220 24480 0 0 $X=256030 $Y=24240
X560 1 155 ICV_15 $T=274620 13600 1 0 $X=274430 $Y=10640
X561 1 7 ICV_15 $T=284280 19040 0 0 $X=284090 $Y=18800
X562 1 181 ICV_15 $T=312340 24480 0 0 $X=312150 $Y=24240
X563 1 2 4 ICV_16 $T=11500 19040 1 0 $X=11310 $Y=16080
X564 1 2 5 ICV_16 $T=11500 24480 1 0 $X=11310 $Y=21520
X565 1 2 6 ICV_16 $T=11500 29920 1 0 $X=11310 $Y=26960
X566 1 2 14 ICV_16 $T=27140 24480 0 0 $X=26950 $Y=24240
X567 1 2 38 ICV_16 $T=66240 35360 1 0 $X=66050 $Y=32400
X568 1 2 221 ICV_16 $T=91080 24480 0 0 $X=90890 $Y=24240
X569 1 2 56 ICV_16 $T=96140 29920 0 0 $X=95950 $Y=29680
X570 1 2 44 ICV_16 $T=117300 29920 1 0 $X=117110 $Y=26960
X571 1 2 81 ICV_16 $T=139380 19040 0 0 $X=139190 $Y=18800
X572 1 2 7 ICV_16 $T=149500 13600 1 0 $X=149310 $Y=10640
X573 1 2 92 ICV_16 $T=160540 29920 0 0 $X=160350 $Y=29680
X574 1 2 96 ICV_16 $T=164220 13600 0 0 $X=164030 $Y=13360
X575 1 2 100 ICV_16 $T=178020 13600 1 0 $X=177830 $Y=10640
X576 1 2 7 ICV_16 $T=179400 19040 1 0 $X=179210 $Y=16080
X577 1 2 103 ICV_16 $T=179860 24480 1 0 $X=179670 $Y=21520
X578 1 2 108 ICV_16 $T=194580 24480 0 0 $X=194390 $Y=24240
X579 1 2 126 ICV_16 $T=217580 19040 1 0 $X=217390 $Y=16080
X580 1 2 9 ICV_16 $T=222640 35360 1 0 $X=222450 $Y=32400
X581 1 2 7 ICV_16 $T=234600 24480 0 0 $X=234410 $Y=24240
X582 1 2 133 ICV_16 $T=236440 29920 1 0 $X=236250 $Y=26960
X583 1 2 134 ICV_16 $T=237360 35360 1 0 $X=237170 $Y=32400
X584 1 2 229 ICV_16 $T=247940 29920 0 0 $X=247750 $Y=29680
X585 1 2 7 ICV_16 $T=262660 29920 1 0 $X=262470 $Y=26960
X586 1 2 7 ICV_16 $T=264960 13600 1 0 $X=264770 $Y=10640
X587 1 2 149 ICV_16 $T=264960 19040 1 0 $X=264770 $Y=16080
X588 1 2 157 ICV_16 $T=277380 19040 0 0 $X=277190 $Y=18800
X589 1 2 7 ICV_16 $T=296700 13600 1 0 $X=296510 $Y=10640
X590 1 2 173 ICV_16 $T=299460 19040 0 0 $X=299270 $Y=18800
X591 1 2 7 ICV_16 $T=306360 13600 1 0 $X=306170 $Y=10640
X592 1 2 182 ICV_16 $T=313260 35360 1 0 $X=313070 $Y=32400
X593 1 2 7 ICV_16 $T=319700 35360 1 0 $X=319510 $Y=32400
X594 1 2 7 ICV_16 $T=320160 19040 1 0 $X=319970 $Y=16080
X595 1 2 186 ICV_16 $T=320620 13600 1 0 $X=320430 $Y=10640
X596 1 2 3 ICV_16 $T=332580 24480 0 0 $X=332390 $Y=24240
X597 1 2 49 2 53 1 sky130_fd_sc_hd__inv_8 $T=91080 29920 0 0 $X=90890 $Y=29680
X598 1 2 56 2 55 1 sky130_fd_sc_hd__inv_8 $T=93840 35360 1 0 $X=93650 $Y=32400
X599 1 2 68 2 71 1 sky130_fd_sc_hd__inv_8 $T=119140 29920 0 0 $X=118950 $Y=29680
X600 1 2 73 2 70 1 sky130_fd_sc_hd__inv_8 $T=122360 35360 1 0 $X=122170 $Y=32400
X601 1 2 79 2 80 1 sky130_fd_sc_hd__inv_8 $T=136160 29920 0 0 $X=135970 $Y=29680
X602 1 2 92 2 95 1 sky130_fd_sc_hd__inv_8 $T=161460 35360 1 0 $X=161270 $Y=32400
X603 1 2 224 2 111 1 sky130_fd_sc_hd__inv_8 $T=189520 24480 1 0 $X=189330 $Y=21520
X604 1 2 228 2 119 1 sky130_fd_sc_hd__inv_8 $T=208380 29920 1 0 $X=208190 $Y=26960
X605 1 2 125 2 127 1 sky130_fd_sc_hd__inv_8 $T=217580 35360 1 0 $X=217390 $Y=32400
X606 1 2 229 2 140 1 sky130_fd_sc_hd__inv_8 $T=245640 35360 1 0 $X=245450 $Y=32400
X607 1 2 158 2 154 1 sky130_fd_sc_hd__inv_8 $T=272780 24480 0 0 $X=272590 $Y=24240
X608 1 2 3 3 9 13 7 ICV_17 $T=7820 13600 0 0 $X=7630 $Y=13360
X609 1 2 3 3 21 27 7 ICV_17 $T=34960 13600 0 0 $X=34770 $Y=13360
X610 1 2 3 3 26 31 7 ICV_17 $T=44160 29920 0 0 $X=43970 $Y=29680
X611 1 2 3 3 42 47 7 ICV_17 $T=70380 19040 0 0 $X=70190 $Y=18800
X612 1 2 3 3 59 64 7 ICV_17 $T=99360 24480 0 0 $X=99170 $Y=24240
X613 1 2 3 3 72 77 7 ICV_17 $T=120060 19040 0 0 $X=119870 $Y=18800
X614 1 2 7 242 223 79 7 ICV_17 $T=128340 24480 0 0 $X=128150 $Y=24240
X615 1 2 78 3 81 85 7 ICV_17 $T=133860 24480 1 0 $X=133670 $Y=21520
X616 1 2 84 3 84 89 7 ICV_17 $T=143980 19040 1 0 $X=143790 $Y=16080
X617 1 2 3 3 88 94 7 ICV_17 $T=147200 19040 0 0 $X=147010 $Y=18800
X618 1 2 3 3 100 105 7 ICV_17 $T=175260 13600 0 0 $X=175070 $Y=13360
X619 1 2 3 3 103 106 7 ICV_17 $T=177560 19040 0 0 $X=177370 $Y=18800
X620 1 2 7 243 225 224 7 ICV_17 $T=180780 29920 0 0 $X=180590 $Y=29680
X621 1 2 130 3 130 135 7 ICV_17 $T=226780 24480 1 0 $X=226590 $Y=21520
X622 1 2 7 3 131 136 7 ICV_17 $T=228160 19040 1 0 $X=227970 $Y=16080
X623 1 2 3 3 132 139 7 ICV_17 $T=232760 19040 0 0 $X=232570 $Y=18800
X624 1 2 7 244 133 229 7 ICV_17 $T=234600 29920 0 0 $X=234410 $Y=29680
X625 1 2 145 3 143 150 7 ICV_17 $T=255300 24480 1 0 $X=255110 $Y=21520
X626 1 2 3 3 149 156 7 ICV_17 $T=263120 13600 0 0 $X=262930 $Y=13360
X627 1 2 3 3 170 176 7 ICV_17 $T=294860 13600 0 0 $X=294670 $Y=13360
X628 1 2 3 3 169 179 7 ICV_17 $T=298080 29920 0 0 $X=297890 $Y=29680
X629 1 2 230 3 177 184 7 ICV_17 $T=304060 24480 1 0 $X=303870 $Y=21520
X630 1 2 3 3 186 191 7 ICV_17 $T=318320 13600 0 0 $X=318130 $Y=13360
X631 1 2 3 3 187 192 7 ICV_17 $T=319240 24480 0 0 $X=319050 $Y=24240
X632 1 2 193 3 194 198 7 ICV_17 $T=332580 19040 1 0 $X=332390 $Y=16080
X633 1 2 44 45 2 220 1 sky130_fd_sc_hd__nor2_4 $T=77280 35360 1 0 $X=77090 $Y=32400
X634 1 2 44 50 2 221 1 sky130_fd_sc_hd__nor2_4 $T=84180 35360 1 0 $X=83990 $Y=32400
X635 1 2 44 63 2 222 1 sky130_fd_sc_hd__nor2_4 $T=109940 29920 0 0 $X=109750 $Y=29680
X636 1 2 44 65 2 69 1 sky130_fd_sc_hd__nor2_4 $T=113620 35360 1 0 $X=113430 $Y=32400
X637 1 2 74 75 2 223 1 sky130_fd_sc_hd__nor2_4 $T=126040 29920 0 0 $X=125850 $Y=29680
X638 1 2 109 110 2 225 1 sky130_fd_sc_hd__nor2_4 $T=189520 35360 1 0 $X=189330 $Y=32400
X639 1 2 109 118 2 226 1 sky130_fd_sc_hd__nor2_4 $T=202860 35360 1 0 $X=202670 $Y=32400
X640 1 2 109 114 2 227 1 sky130_fd_sc_hd__nor2_4 $T=203320 29920 0 0 $X=203130 $Y=29680
X641 1 2 173 230 2 1 sky130_fd_sc_hd__clkbuf_1 $T=301760 24480 1 0 $X=301570 $Y=21520
X642 1 2 230 2 174 1 sky130_fd_sc_hd__clkbuf_4 $T=301760 29920 1 0 $X=301570 $Y=26960
X643 1 2 155 2 164 1 sky130_fd_sc_hd__clkbuf_16 $T=277840 13600 1 0 $X=277650 $Y=10640
X644 1 2 3 5 11 7 ICV_41 $T=7820 24480 0 0 $X=7630 $Y=24240
X645 1 2 3 16 23 7 ICV_41 $T=33580 24480 1 0 $X=33390 $Y=21520
X646 1 2 3 33 40 7 ICV_41 $T=61640 29920 1 0 $X=61450 $Y=26960
X647 1 2 3 48 57 7 ICV_41 $T=88780 19040 1 0 $X=88590 $Y=16080
X648 1 2 3 96 99 7 ICV_41 $T=161460 19040 1 0 $X=161270 $Y=16080
X649 1 2 3 117 123 7 ICV_41 $T=201940 19040 1 0 $X=201750 $Y=16080
X650 1 2 245 124 9 7 ICV_41 $T=215740 29920 0 0 $X=215550 $Y=29680
X651 1 2 3 138 142 7 ICV_41 $T=243800 13600 0 0 $X=243610 $Y=13360
X652 1 2 3 157 162 7 ICV_41 $T=273700 24480 1 0 $X=273510 $Y=21520
X653 1 2 3 160 166 7 ICV_41 $T=281520 19040 1 0 $X=281330 $Y=16080
X654 1 2 3 161 167 7 ICV_41 $T=282440 35360 1 0 $X=282250 $Y=32400
X655 1 2 3 168 178 7 ICV_41 $T=297160 24480 0 0 $X=296970 $Y=24240
X656 1 2 3 175 183 7 ICV_41 $T=304520 19040 1 0 $X=304330 $Y=16080
X657 1 2 3 181 188 7 ICV_41 $T=314180 29920 1 0 $X=313990 $Y=26960
X658 1 2 3 185 190 7 ICV_41 $T=319700 29920 0 0 $X=319510 $Y=29680
X659 1 2 3 195 199 7 ICV_41 $T=334420 35360 1 0 $X=334230 $Y=32400
X660 1 2 3 193 200 7 ICV_41 $T=334880 24480 1 0 $X=334690 $Y=21520
.ENDS
***************************************
.SUBCKT deserialiser_unit_cell_1 VSS VDD PAR_IN4<29> OUT<7> OUT<2> PAR_IN2<10> COMPLETE PAR_IN5<29> PAR_IN2<22> RESET PAR_IN6<15> PAR_IN7<22> PAR_IN7<7> PAR_IN6<14> OUT<9> PAR_IN8<19> PAR_IN1<14> PAR_IN1<1> PAR_IN4<8> PAR_IN4<12>
+ INTERNAL_FINISH PAR_IN6<13> OUT<6> PAR_IN8<3> PAR_IN8<5> COUNT<4> OUT<10> OUT<26> OUT<11> PAR_IN3<12> PAR_IN7<6> PAR_IN6<22> PAR_IN1<25> OUT<22> OUT<23> PAR_IN8<28> PAR_IN8<13> PAR_IN3<25> PAR_IN1<30> OUT<15>
+ PAR_IN2<8> OUT<25> OUT<16> PAR_IN5<7> READY PAR_IN2<9> PAR_IN4<25> PAR_IN4<3> PAR_IN7<13> PAR_IN8<14> PAR_IN5<1> PAR_IN2<5> PAR_IN6<8> PAR_IN5<21> PAR_IN3<19> PAR_IN6<4> PAR_IN2<4> OUT<0> PAR_IN5<19> PAR_IN1<24>
+ PAR_IN3<26> PAR_IN1<12> PAR_IN6<23> PAR_IN4<20> PAR_IN4<22> PAR_IN8<31> PAR_IN4<0> PAR_IN5<12> PAR_IN7<9> PAR_IN5<9> COUNT<3> PAR_IN7<1> PAR_IN2<19> PAR_IN3<1> PAR_IN8<9> PAR_IN8<26> PAR_IN6<28> PAR_IN4<14> PAR_IN3<24> PAR_IN5<5>
+ PAR_IN7<25> PAR_IN6<7> PAR_IN7<3> PAR_IN5<18> PAR_IN8<20> PAR_IN4<23> PAR_IN1<26> PAR_IN7<19> PAR_IN3<31> PAR_IN6<25> PAR_IN3<0> PAR_IN7<0> PAR_IN1<8> PAR_IN6<10> PAR_IN5<4> OUT<13> PAR_IN6<29> PAR_IN6<6> PAR_IN5<14> PAR_IN5<13>
+ PAR_IN4<10> PAR_IN5<0> PAR_IN7<8> PAR_IN4<13> PAR_IN5<6> SAMPLE_COUNT<2> PAR_IN7<5> PAR_IN6<12> PAR_IN5<17> SAMPLE_COUNT<1> COUNT<1> PAR_IN2<28> PAR_IN5<20> PAR_IN4<15> PAR_IN8<2> OUT<5> PAR_IN3<14> PAR_IN8<10> PAR_IN4<5> OUT<4>
+ OUT<1> PAR_IN8<25> OUT<28> PAR_IN2<18> OUT<24> COUNT<2> COUNT<0> PAR_IN3<3> PAR_IN8<24> PAR_IN5<11> PAR_IN7<4> PAR_IN6<19> PAR_IN4<4> PAR_IN6<16> OUT<3> PAR_IN3<8> PAR_IN3<29> OUT<12> PAR_IN5<15> OUT<18>
+ OUT<21> OUT<17> COUNT<5> OUT<30> OUT<31> SAMPLE_COUNT<3> SAMPLE_COUNT<0> PAR_IN3<22> PAR_IN1<3> PAR_IN5<25> PAR_IN3<20> PAR_IN2<1> PAR_IN5<16> PAR_IN5<8> PAR_IN6<30> PAR_IN7<21> PAR_IN5<28> PAR_IN4<21> PAR_IN4<27> PAR_IN8<17>
+ PAR_IN2<20> PAR_IN2<31> PAR_IN2<24> PAR_IN5<27> PAR_IN7<20> PAR_IN7<23> PAR_IN1<16> OUT<19> PAR_IN1<31> PAR_IN3<5> PAR_IN7<10> PAR_IN8<4> PAR_IN7<17> PAR_IN1<11> OUT<14> PAR_IN2<29> PAR_IN2<11> PAR_IN5<10> PAR_IN2<30> OUT<20>
+ PAR_IN7<14> PAR_IN1<21> PAR_IN2<25> PAR_IN4<19> PAR_IN2<14> PAR_IN3<15> PAR_IN4<18> PAR_IN8<8> CLK PAR_IN1<13> PAR_IN7<31> PAR_IN1<4> PAR_IN4<6> PAR_IN5<22> PAR_IN7<24> PAR_IN8<12> OUT<29> PAR_IN3<6> PAR_IN8<29> PAR_IN4<9>
+ PAR_IN4<31> PAR_IN3<28> PAR_IN6<1> PAR_IN2<2> PAR_IN6<21> PAR_IN8<1> PAR_IN7<11> SERIAL_IN PAR_IN3<27> PAR_IN8<11> PAR_IN4<16> PAR_IN8<18> PAR_IN4<1> PAR_IN1<17> PAR_IN2<6> PAR_IN6<17> OUT<27> PAR_IN6<20> PAR_IN7<18> PAR_IN2<0>
+ PAR_IN3<18> PAR_IN8<15> PAR_IN7<27> PAR_IN5<30> PAR_IN6<26> PAR_IN1<9> PAR_IN8<30> PAR_IN4<11> PAR_IN3<4> PAR_IN2<17> PAR_IN4<17> PAR_IN8<0> PAR_IN6<9> PAR_IN2<26> PAR_IN1<0> PAR_IN6<3> PAR_IN3<30> PAR_IN8<16> PAR_IN6<24> PAR_IN3<9>
+ PAR_IN7<2> PAR_IN1<20> PAR_IN1<28> PAR_IN2<27> PAR_IN7<16> PAR_IN7<12> PAR_IN1<5> PAR_IN4<24> PAR_IN6<11> PAR_IN6<5> PAR_IN3<23> PAR_IN6<27> PAR_IN5<23> PAR_IN6<18> PAR_IN8<21> PAR_IN2<13> PAR_IN8<27> PAR_IN4<2> PAR_IN1<7> PAR_IN8<22>
+ PAR_IN1<15> PAR_IN2<16> PAR_IN6<0> PAR_IN1<22> PAR_IN3<21> PAR_IN8<23> PAR_IN5<26> PAR_IN2<7> PAR_IN2<12> PAR_IN7<15> PAR_IN2<15> PAR_IN1<27> PAR_IN4<26> PAR_IN1<10> PAR_IN7<26> PAR_IN7<28> PAR_IN3<11> PAR_IN1<2> PAR_IN1<19> PAR_IN3<7>
+ OUT<8> PAR_IN1<18> PAR_IN1<6> PAR_IN2<21> PAR_IN3<2> PAR_IN8<7> PAR_IN7<30> PAR_IN1<23> PAR_IN8<6> PAR_IN3<13> PAR_IN5<2> PAR_IN2<3> PAR_IN4<7> PAR_IN3<10> PAR_IN5<3> PAR_IN4<28> PAR_IN5<31> PAR_IN3<17> PAR_IN1<29> PAR_IN5<24>
+ PAR_IN3<16> PAR_IN2<23> PAR_IN6<31> PAR_IN6<2> PAR_IN7<29> PAR_IN4<30>
** N=1116 EP=306 IP=2857 FDC=63394
X0 VSS VDD Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=123705 $D=191
X1 VSS VDD Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=172665 $D=191
X2 VSS VDD Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=216185 $D=191
X3 VSS VDD Dpar a=977.425 p=696.42 m=1 $[nwdiode] $X=5330 $Y=308665 $D=191
X4 1115 VDD Probe probetype=1 $[VDD] $X=178018 $Y=27288 $D=314
X5 1116 VSS Probe probetype=1 $[VSS] $X=178018 $Y=103878 $D=314
X6 VSS VDD COMPLETE RESET 19 11 8 12 100 9 16 PAR_IN6<26> PAR_IN8<30> PAR_IN3<4> PAR_IN2<17> PAR_IN8<0> PAR_IN2<10> 20 163 18
+ PAR_IN5<29> 60 50 185 PAR_IN1<9> PAR_IN4<11> PAR_IN6<15> PAR_IN4<17> PAR_IN4<29> PAR_IN2<22> 25 PAR_IN7<22> 139 24 26 PAR_IN7<7> 34 28 32 31
+ PAR_IN6<14> PAR_IN8<19> 68 33 72 41 40 PAR_IN4<8> PAR_IN4<12> 30 45 44 39 PAR_IN1<1> PAR_IN1<14> 37 52 53 PAR_IN2<5> 49
+ PAR_IN2<8> 47 PAR_IN2<9> 55 59 PAR_IN6<13> PAR_IN3<12> 56 144 64 PAR_IN8<3> 67 PAR_IN8<5> PAR_IN7<6> 54 71 73 76 69 PAR_IN2<19>
+ PAR_IN6<22> 87 81 PAR_IN1<12> 79 159 98 82 83 85 88 86 90 PAR_IN5<12> PAR_IN1<25> 95 PAR_IN8<28> PAR_IN7<9> 106 184
+ 93 113 96 99 92 PAR_IN3<25> PAR_IN8<13> 116 107 PAR_IN4<3> 111 109 108 103 112 PAR_IN5<7> 117 114 120 PAR_IN7<1>
+ PAR_IN4<0> PAR_IN7<13> 123 PAR_IN4<25> 124 130 43 126 140 129 127 133 PAR_IN2<4> PAR_IN5<1> 132 134 PAR_IN5<9> 143 137 141
+ PAR_IN3<19> 150 PAR_IN6<4> 153 166 146 PAR_IN5<19> 155 148 152 154 PAR_IN1<30> 156 158 165 PAR_IN1<24> 181 161 171 164
+ PAR_IN6<8> 176 169 PAR_IN3<26> 183 175 173 172 178 PAR_IN4<20> PAR_IN8<14> PAR_IN4<22> 179 186 177 191 188 200 PAR_IN8<9> 199
+ 193 189 195 PAR_IN3<1> PAR_IN8<26> 204 206 202 201 PAR_IN4<14> 207 210 PAR_IN3<24> PAR_IN6<7> PAR_IN5<5> PAR_IN8<31> PAR_IN6<28> 211 213 215
+ 149 216 218 PAR_IN7<3> 212 220 PAR_IN5<18> 226 PAR_IN6<23> 222 197 224 227 232 PAR_IN4<23> 230 229 221 PAR_IN7<25> 228
+ 233 237 PAR_IN1<26> 236 PAR_IN5<21> 238 240 234 PAR_IN7<19> 242 PAR_IN8<16> 243 PAR_IN8<20> 75 PAR_IN3<31> 246 PAR_IN6<25> PAR_IN7<0> 245 196
+ 36 PAR_IN1<8> PAR_IN1<0> PAR_IN6<10> PAR_IN6<3> PAR_IN6<9> PAR_IN2<26> PAR_IN3<30> PAR_IN3<9> PAR_IN6<24> PAR_IN5<4>
+ ICV_20 $T=0 0 0 0 $X=0 $Y=309800
X7 VSS VDD COMPLETE 258 RESET 259 161 343 284 260 PAR_IN1<28> PAR_IN7<2> PAR_IN6<29> PAR_IN1<5> PAR_IN6<6> PAR_IN7<16> PAR_IN7<12> PAR_IN5<14> 263 33
+ PAR_IN1<20> 262 20 PAR_IN5<13> PAR_IN2<27> PAR_IN5<0> PAR_IN7<8> PAR_IN4<10> 24 PAR_IN4<13> 268 270 26 28 25 269 31 34 32 37
+ 40 271 278 177 44 294 273 189 275 52 49 56 55 272 287 53 307 193 54 274
+ 276 295 83 283 279 64 72 280 73 282 76 285 286 281 289 293 79 86 329 290
+ 137 90 288 291 88 82 87 85 292 92 296 297 95 96 113 99 299 302 108 301
+ 303 300 11 112 117 114 109 111 16 304 313 116 305 312 129 107 342 317 298 308
+ 311 314 310 126 123 124 133 309 127 315 322 132 318 321 134 316 319 140 320 141
+ 324 155 148 323 277 337 152 150 325 149 154 334 98 156 158 331 330 327 164 328
+ 93 336 332 333 166 181 171 345 340 172 188 176 178 338 183 339 306 173 191 326
+ 195 200 163 199 341 351 202 344 204 355 206 216 347 346 348 350 211 230 210 354
+ 335 352 353 213 215 349 218 19 220 224 357 227 358 356 359 229 363 360 368 226
+ 233 361 228 236 362 366 242 364 232 240 367 243 369 365 130 81 370 371 PAR_IN3<23> PAR_IN5<6>
+ PAR_IN3<0> PAR_IN6<12> PAR_IN6<18> PAR_IN6<11> PAR_IN6<27> PAR_IN7<5> PAR_IN6<5> PAR_IN4<24> PAR_IN5<23>
+ ICV_25 $T=0 0 0 0 $X=0 $Y=263600
X8 VSS VDD COMPLETE RESET 394 377 282 PAR_IN8<21> PAR_IN2<13> PAR_IN8<27> PAR_IN1<7> PAR_IN5<17> 378 380 398 262 379 PAR_IN4<2> 381 20
+ 9 383 404 389 382 386 384 390 268 387 385 388 269 393 396 45 39 37 395 270
+ 272 271 392 52 24 294 75 391 400 273 278 54 189 274 399 275 401 411 402 41
+ 407 276 403 405 397 406 408 410 279 69 409 280 193 416 71 177 284 53 449 412
+ 413 288 286 285 291 283 292 414 293 59 79 296 289 418 297 85 417 93 419 423
+ 420 421 95 422 424 100 426 103 302 427 428 430 429 425 432 16 431 303 304 305
+ 129 361 331 433 312 349 328 335 326 434 482 311 436 442 435 440 479 362 437 314
+ 322 316 438 448 320 295 444 319 18 315 445 323 443 446 318 321 447 441 450 452
+ 332 324 454 455 325 144 451 83 453 327 330 329 333 460 338 456 458 459 485 461
+ 457 462 179 439 464 339 169 465 463 173 175 360 466 184 467 356 468 358 366 469
+ 344 368 476 471 470 472 473 474 346 370 139 347 353 212 475 351 477 352 481 480
+ 348 355 484 483 486 221 491 359 357 488 492 364 363 489 238 490 493 487 232 495
+ 496 500 498 371 345 499 478 497 PAR_IN8<22> PAR_IN1<15> PAR_IN2<16> PAR_IN5<20> PAR_IN1<22> PAR_IN6<0>
+ ICV_31 $T=0 0 0 0 $X=0 $Y=217360
X9 VSS VDD COMPLETE RESET 403 377 PAR_IN4<15> PAR_IN8<2> PAR_IN8<23> PAR_IN2<7> PAR_IN2<12> PAR_IN5<26> 505 508 259 378 387 506 381 384
+ 507 380 382 388 389 385 383 515 379 391 511 510 521 512 390 30 392 513 509 517
+ 393 516 514 395 394 43 400 83 56 562 405 558 401 177 397 518 398 12 406 519
+ 402 404 520 527 524 407 523 522 532 607 408 67 411 409 525 535 526 531 528 529
+ 556 410 553 530 478 533 534 499 260 414 536 537 95 422 421 418 419 538 541 420
+ 290 539 263 540 544 137 299 427 545 428 424 542 546 547 543 584 245 93 431 426
+ 430 432 550 548 549 551 68 552 555 563 554 436 60 557 328 120 439 437 565 362
+ 561 335 361 560 564 314 438 440 567 566 443 442 441 349 307 315 446 568 308 447
+ 445 444 559 323 320 570 576 293 573 153 589 569 448 585 571 574 453 455 575 452
+ 577 461 456 52 454 459 578 159 460 258 582 579 583 37 458 581 580 596 587 594
+ 588 464 465 590 586 592 466 593 278 467 294 197 469 468 595 608 598 471 473 600
+ 470 472 572 334 597 481 474 343 477 599 476 480 602 449 483 475 336 79 85 601
+ 484 603 358 462 485 492 237 488 493 450 222 491 489 604 490 368 605 496 495 366
+ 606 279 500 PAR_IN8<10> PAR_IN4<5> PAR_IN7<15> PAR_IN2<28> PAR_IN1<27> PAR_IN2<15>
+ ICV_33 $T=0 0 0 0 $X=0 $Y=173800
X10 VSS VDD COMPLETE RESET 614 451 381 PAR_IN3<21> PAR_IN8<25> 380 505 615 645 507 509 508 506 512 617 511
+ 619 621 618 513 537 540 515 514 517 43 516 47 519 520 521 620 50 524 527 626
+ 624 559 622 523 522 525 526 625 568 623 529 531 631 532 530 629 630 533 534 632
+ 634 536 633 628 627 535 654 543 635 539 638 542 593 641 545 547 639 544 637 546
+ 640 550 642 560 571 549 579 555 643 557 552 644 548 570 299 646 558 246 561 647
+ 328 650 361 335 562 563 564 648 565 349 649 290 566 651 652 567 326 653 362 573
+ 574 146 661 159 590 577 636 656 578 581 580 657 582 165 655 584 583 658 585 592
+ 588 659 594 662 660 595 360 497 358 356 366 663 368 599 668 664 666 185 671 670
+ 667 665 669 600 426 336 673 672 674 602 678 604 222 679 675 677 676 682 681 680
+ 683 607 608 PAR_IN4<26> PAR_IN7<26> PAR_IN1<10>
+ ICV_34 $T=0 0 0 0 $X=0 $Y=149360
X11 VSS VDD COMPLETE RESET PAR_IN7<28> PAR_IN3<11> 684 708 710 560 686 687 385 392 688 689 386 36 618 648
+ 391 400 47 690 691 715 753 693 695 519 694 692 622 OUT<10> 624 685 627 628 626 696
+ 697 629 699 698 OUT<22> OUT<23> OUT<26> 630 700 703 631 702 633 541 701 632 635 705 636 660
+ 637 638 OUT<25> 706 546 653 639 707 545 641 712 711 709 540 557 713 505 644 716 645
+ 313 299 646 649 714 647 717 754 650 651 514 718 287 324 307 652 654 326 734 143
+ 719 720 722 721 737 724 106 735 723 733 726 727 728 729 655 165 730 731 725 732
+ 570 196 736 186 738 201 661 741 739 614 740 662 663 742 745 599 743 744 666 665
+ 670 746 669 668 667 602 365 368 747 748 672 671 79 673 674 85 679 677 678 676
+ 334 749 675 335 750 681 752 751 683 682 680 634 PAR_IN1<2> PAR_IN3<14> PAR_IN3<7> PAR_IN1<19>
+ ICV_35 $T=0 0 0 0 $X=0 $Y=124880
X12 VSS VDD 317 840 828 838 836 872 843 827 COMPLETE RESET 620 623 615 685 686 PAR_IN2<18> PAR_IN1<18> PAR_IN1<6>
+ PAR_IN2<21> 756 8 687 688 757 758 389 759 560 509 689 512 540 732 711 OUT<7> OUT<8> 396 731
+ 761 648 765 764 OUT<9> 766 763 762 537 690 691 767 OUT<13> OUT<6> 770 693 769 773 695 772
+ 775 771 391 768 774 694 776 OUT<10> 777 779 OUT<11> 780 789 400 782 698 783 784 696 OUT<24>
+ 625 697 787 700 785 OUT<22> 791 786 788 790 699 702 792 706 703 794 778 793 801 798
+ 797 795 799 796 705 636 817 800 811 OUT<28> 810 816 803 805 809 593 804 806 807 579
+ 707 814 815 808 812 709 813 COUNT<2> 571 COUNT<0> COUNT<1> 802 643 COUNT<3> 710 818 819 708 826 713
+ 823 821 313 397 845 822 837 READY 714 841 831 824 829 833 825 832 OUT<0> 715 835 834
+ 650 293 718 846 441 287 736 569 723 324 720 844 839 568 307 847 842 721 719 848
+ 849 514 850 725 726 724 727 851 728 735 878 656 729 589 730 733 737 853 485 432
+ 861 443 639 852 462 860 862 738 855 657 859 641 854 856 585 858 857 740 863 871
+ 866 SAMPLE_COUNT<1> 627 864 760 741 SAMPLE_COUNT<2> 865 739 868 742 869 870 660 867 745 876 874 746 479
+ 873 350 365 875 880 877 482 674 354 748 879 734 649 299 881 882 883 234 884 887
+ 886 885 891 369 890 888 889 749 893 892 750 753 337 663 587 596 342 606 PAR_IN3<2> PAR_IN3<13>
+ 754 PAR_IN1<23> PAR_IN3<3> PAR_IN8<7> PAR_IN8<6> PAR_IN7<30> PAR_IN5<2> PAR_IN5<11> PAR_IN8<24>
+ ICV_38 $T=0 0 0 0 $X=0 $Y=78640
X13 VSS VDD COUNT<4> 835 834 847 COMPLETE RESET 684 281 309 554 347 620 617 PAR_IN7<4> PAR_IN3<10> PAR_IN5<3> PAR_IN4<28> PAR_IN5<31>
+ PAR_IN6<19> 756 341 269 PAR_IN2<3> 757 412 OUT<4> 851 PAR_IN6<16> PAR_IN4<7> 759 OUT<2> OUT<1> PAR_IN3<8> 762 OUT<3> 763 767 PAR_IN3<29>
+ PAR_IN4<4> 766 OUT<5> 761 765 298 764 772 823 OUT<12> 769 PAR_IN5<15> 774 768 909 771 777 773 906 907
+ 815 770 OUT<18> 913 807 775 911 776 779 784 804 780 778 910 786 912 782 790 568 627
+ 783 559 628 787 OUT<21> 806 785 788 792 916 915 789 397 919 791 OUT<15> 917 808 793 918
+ 794 532 920 553 797 798 556 795 813 OUT<17> OUT<16> 800 812 802 799 805 803 810 922 INTERNAL_FINISH
+ 811 818 COUNT<5> 809 924 OUT<30> 814 824 826 COUNT<2> 816 941 817 READY 926 819 822 821 570 825
+ 832 827 927 OUT<31> 828 649 829 836 831 443 833 840 930 837 929 839 864 934 848 842
+ 931 838 841 933 843 935 932 845 844 846 936 574 726 937 619 COUNT<0> 889 621 939 850
+ 299 940 432 942 943 853 658 884 854 944 855 SAMPLE_COUNT<3> 858 863 945 SAMPLE_COUNT<0> 859 869 856 860
+ 861 656 589 865 947 SAMPLE_COUNT<2> 948 862 SAMPLE_COUNT<1> 875 641 950 866 867 868 872 870 207 871 873
+ 881 485 876 874 877 951 878 674 879 880 885 PAR_IN3<22> 883 952 954 882 955 956 886 887
+ 890 888 892 891 893 938 659 709 717 498 PAR_IN3<17> PAR_IN1<29> PAR_IN2<23> PAR_IN1<3> PAR_IN3<16> PAR_IN5<24> PAR_IN6<31>
+ ICV_40 $T=0 0 0 0 $X=0 $Y=35120
X14 VSS VDD COMPLETE 433 760 277 RESET 347 939 PAR_IN5<25> PAR_IN3<20> PAR_IN6<2> PAR_IN2<1> 310 301 743 758 PAR_IN5<16> 306 PAR_IN5<8>
+ 425 510 PAR_IN7<21> PAR_IN3<5> PAR_IN6<30> 463 PAR_IN5<28> PAR_IN2<11> 564 572 PAR_IN4<21> 518 945 906 PAR_IN4<27> 692 PAR_IN8<17> 907 PAR_IN2<14> PAR_IN2<31>
+ PAR_IN2<20> 701 OUT<18> 909 910 429 PAR_IN2<24> 664 OUT<19> 912 744 PAR_IN5<27> 911 528 913 OUT<20> PAR_IN7<20> PAR_IN1<16> 409 PAR_IN7<23>
+ 413 915 917 PAR_IN1<11> 918 538 PAR_IN7<10> OUT<14> 920 919 916 597 OUT<17> 794 796 PAR_IN8<4> PAR_IN7<17> 300 OUT<27> 801
+ 640 924 635 642 PAR_IN2<29> PAR_IN5<10> 922 430 PAR_IN2<30> OUT<30> PAR_IN1<21> OUT<29> 926 PAR_IN7<14> 802 712 435 927 PAR_IN2<25> 438
+ PAR_IN4<19> OUT<31> 416 839 PAR_IN4<18> PAR_IN1<13> PAR_IN3<15> 716 841 929 930 842 931 932 274 PAR_IN1<4> 575 933 936 PAR_IN4<6>
+ 935 399 PAR_IN8<8> 937 938 759 934 PAR_IN4<9> PAR_IN3<6> 849 457 586 942 943 PAR_IN4<31> PAR_IN8<29> 340 852 PAR_IN8<12> 940
+ PAR_IN3<28> 551 PAR_IN6<1> 948 947 417 PAR_IN2<2> 857 PAR_IN8<1> 950 PAR_IN1<31> PAR_IN7<11> 941 CLK PAR_IN3<27> 598 SERIAL_IN 576 359 951
+ PAR_IN8<11> PAR_IN4<16> 952 747 PAR_IN6<21> PAR_IN7<31> 630 513 601 423 PAR_IN7<24> 955 954 487 PAR_IN8<18> 486 PAR_IN1<17> PAR_IN2<6> PAR_IN4<1> 944
+ 956 PAR_IN5<22> PAR_IN6<17> 367 603 605 PAR_IN2<0> 751 PAR_IN6<20> PAR_IN8<15> PAR_IN7<18> 752 434 722 PAR_IN7<27> PAR_IN3<18> PAR_IN5<30> PAR_IN4<30> PAR_IN7<29>
+ ICV_42 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
